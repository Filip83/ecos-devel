#==========================================================================
#
#       kbd_button.cdl
#
#       eCos configuration data for the Atmel AVR32 button keyboard driver
#
#==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
#==========================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    Filip
# Contributors:
# Date:         2016-11-23
# Purpose:
# Description:  Button keyboard driver for Atmel AVR32
#
#####DESCRIPTIONEND####
#
#==========================================================================

cdl_package CYGPKG_DEVS_KBD_BUTTON {
    display     "Button keyboard driver."
    include_dir cyg/io

    active_if   CYGPKG_IO_FILEIO
    requires    CYGPKG_IO
    requires    CYGFUN_KERNEL_API_C

    compile       -library=libextras.a kbd_matrix.c

    description "Keyboard driver for the button"

    cdl_component CYGPKG_DEVS_KBD_BUTTON_OPTIONS {
        display "options"
        flavor  none
        no_define

        cdl_option CYGPKG_DEVS_KBD_BUTTON_CFLAGS {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description "
               This option modifies the set of compiler flags for
               building the keypad driver package. These flags
               are used in addition to the set of global flags."
        }

        cdl_option CYGDAT_DEVS_KBD_BUTTON_NAME {
            display "Device name for the keyboard driver"
            flavor data
            default_value {"\"/dev/kbd\""}
            description " This option specifies the name of the keypad device"
        }

        cdl_option CYGNUM_DEVS_KBD_BUTTON_SCAN_INTERVAL {
            display "Keyboard scan interval"
            flavor data
            legal_value   1 to 128
            default_value { 7 }
            description "
                This option defines keyboard scan interval.
                This interval is used for glitch filter and key
                repeat scan."
        }

        cdl_option CYGNUM_DEVS_KBD_BUTTON_NUM_IO_INTERRUPTS_GROUP {
            display "Numer to gpio interrupst gorups to use"
            flavor data
            legal_value   1 to 4
            default_value { 1 }
            description "
                This option defines nuber of gpio interrupt groups.
                The value of this option must be set to number of
                interrupt group to which button are connected."
        }

        cdl_option CYGNUM_DEVS_KBD_MATRIX_BUTTON_MODE {
            display "Keyboard driver callback mode"
            flavor bool
            default_value { 0 }
            description "
                This option enable callback only mode. In this mode
                callback function to deliver key strokes is used.
                Keyboard IO functionality is disabled."
        }

        cdl_option CYGNUM_DEVS_KBD_BUTTON_INTERRUPT_PRIO {
            display "Keyboard driver interrupt priority"
            flavor data
            legal_values  0 to 3
            default_value { 0 }
            description "
                This option set keyboard river insterrupt priortiy."
        }

        cdl_option CYGNUM_DEVS_KBD_BUTTON_EVENT_BUFFER_SIZE {
            display "Number of events the driver can buffer"
            active_if CYGNUM_DEVS_KBD_MATRIX_CALLBACK_MODE == 0
            flavor data
            default_value { 5 }
            description "
                This option defines the size of the keypad device internal
            buffer. The cyg_io_read() function will return as many of these
            as there is space for in the buffer passed."
        }
    }
}
