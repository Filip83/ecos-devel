# ====================================================================
#
#      flash_avr32_uc3c.cdl
#
#      Atmel AVR32UC3C flash memory package
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Contributors:
# Date:           2012-11-15
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_AVR32_CDW {
    display     "AVR32 internal FLASHCDW memory support"
    description "Support for the internal FLASH memory of AVR32UC3C controllers"

    parent      CYGPKG_IO_FLASH
    active_if   CYGPKG_IO_FLASH
    requires    CYGPKG_HAL_AVR32
    implements  CYGHWR_IO_FLASH_DEVICE

    include_dir   cyg/io
    compile -library=libextras.a flash_avr32_cdw.c flashcdw.c
    

    cdl_option CYGPKG_DEVS_FLASH_AVR32_CDW_START {
         display "FLASH region start address"
         flavor  data
         default_value 0x80000000
         description   "
             This option specifies the start address of internal FLASH
             memory to access with this driver."
    }

    cdl_option CYGPKG_DEVS_FLASH_AVR32_CDW_END {
         display "FLASH region end address"
         flavor  data
         default_value 0x80040000
         description   "
             This option specifies the end address of internal FLASH
             memory to access with this driver."
    }

}
