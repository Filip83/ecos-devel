##=============================================================================
##
##      spi_ltc2600.cdl
##
##      LTC2600 SPI dac driver configuration options.
##
##=============================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##=============================================================================
#######DESCRIPTIONBEGIN####
##
##
## Author(s):   Mike Jones
## Date:        2013-06-13
## Purpose:     Configure LTC SPI dac driver.
##
######DESCRIPTIONEND####
##
##=============================================================================

cdl_package CYGPKG_DEVS_DAC_SPI_LTC2600 {
    display      "Linear Technology LTC2600 DAC support"
    parent        CYGPKG_IO_DAC_DEVICES
    active_if     { CYGPKG_IO_DAC_DEVICES && CYGPKG_IO_SPI }
    requires      {CYGNUM_IO_DAC_OUTPUT_SIZE >= 16}
    description "
        This option enables the DAC device drivers for the LTC2600 on the TWR-ADCDAC-LTC"

    include_dir   cyg/io
    compile       -library=libextras.a dac_ltc2600.c

    cdl_interface CYGHWR_DEVS_DAC_SPI_LTC2600_DEVICE {
        display     "Hardware LTC2600 DAC device drivers"
        description "
            This calculated option gives the number of DAC2600 dac
            devices on the current platform."
    }

     cdl_option CYGPKG_DEVS_DAC_LTC2600_TRACE {
        display       "DAC driver tracing"
        flavor        bool
        default_value 0
        description   "
            Enable tracing of the DAC driver. Select to debug the driver."
    }

    cdl_component CYGHWR_DEVS_DAC_LTC2600_DAC1 {
        display         "DAC1"
        default_value   0
        description     "
            DAC1 supports 8 analog output channels."
        
        cdl_interface CYGINT_DEVS_DAC_LTC2600_DAC1_CHANNELS {
            display         "Number of DAC channels"
        }
                    
        cdl_option CYGNUM_DEVS_DAC_LTC2600_DAC1_DEFAULT_RATE {
            display         "Default sample rate"
            flavor          data
            legal_values    1 to 100000
            default_value   1000
            description     "
                The driver will be initialized with the default sample rate.
                If you raise the default sample rate you might need to increase
                the buffer size for each channel."
        }
             
        cdl_option CYGNUM_DEVS_DAC_LTC2600_DAC1_TMR {
            display         "Timer unit"
            flavor          data
            legal_values    0 to 2
            default_value   1
            description     "
                The DAC will use the slected timer
                module to generate interrupts. 0-1 is the FTM
                module and 2 is the PDB module. The choice
                of timer modules affects the achievable sample
                rate. FTM and PDB can divide down the system
                clock with a 16 bit counter. However, the PDB
                also has two prescalers, one that scales from
                a 1X-40X, and one that scales from 1X-128X."
        }
   
        cdl_option CYGNUM_DEVS_DAC_LTC2600_DAC1_TMR_INT_PRI {
            display         "TMR interrupt priority"
            flavor          data
            default_value   0x80
            description     "
                Priority of the timer module request interrupt."
        }

        # DAC1 supports 8 analog outputs
        for { set ::channel 0 } { $::channel < 8 } { incr ::channel } {  
    
            cdl_component CYGHWR_DEVS_DAC_LTC2600_DAC1_CHANNEL[set ::channel] {
                display         "DAC channel [set ::channel]"
                flavor          bool
                default_value   [set ::channel] == 0
                implements      CYGINT_DEVS_DAC_LTC2600_DAC1_CHANNELS
                description     "
                    If the application needs to access the DAC
                    channel [set ::channel] via an eCos DAC driver then
                    this option should be enabled."
     
                cdl_option CYGDAT_DEVS_DAC_LTC2600_DAC1_CHANNEL[set ::channel]_NAME {
                    display         "Device name"
                    flavor          data
                    default_value   [format {"\"/dev/dac1%d\""} $::channel]
                    description     "
                        This option controls the name that an eCos application
                        should use to access this device via cyg_io_lookup(),
                        open(), or similar calls."
                }
        
                cdl_option CYGDAT_DEVS_DAC_LTC2600_DAC1_CHANNEL[set ::channel]_BUFSIZE {
                    display         "Size of data buffer"
                    flavor          data
                    legal_values    1 to 65536
                    default_value   128
                    description     "
                        This option controls the amount of data the
                        buffer can store. The required RAM is = size of
                        data buffer * 2."
                } 
            }
        }
    }
        
    cdl_component CYGPKG_DEVS_DAC_SPI_LTC2600_TESTS {
        display         "LTC2600 tests"
        flavor          data
        active_if       CYGPKG_KERNEL
        active_if       CYGPKG_IO_SPI
        active_if       { CYGHWR_DEVS_DAC_SPI_LTC2600_DEVICE >= 1 }
        no_define
        calculated      { "tests/dac_ltc2600_test.c" }
        description     "
            This option specifies the set of tests for ltc2600 driver."
    }
}

# EOF spi_ltc2600.cdl
