# ====================================================================
#
#      bluetooth.cdl
#
#      Bluetooth stack to implement comunication via bluetooth.
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2003 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip 
# Contributors:   
# Date:           2018-12-16
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_BLUETOOTH_LIB {
    display         "Bletooth stack"
    include_dir     btlib

    requires        CYGPKG_ISOINFRA
    requires        CYGPKG_MEMALLOC
    requires        CYGPKG_ERROR
    
    compile         -library=libextras.a\
    				ad_parser.c \
					ant_cmd.c \
					bluetooth_init_cc2560B_1.4_BT_Spec_4.1.c \
					btstack_chipset_cc256x.c \
					btstack_linked_list.c \
					btstack_memory.c \
					btstack_memory_pool.c \
					btstack_ring_buffer.c \
					btstack_run_loop.c \
					btstack_run_loop_ecos.c \
					btstack_slip.c \
					btstack_util.c \
					hci.c \
					hci_cmd.c \
					hci_dump.c \
					hci_transport_h4.c \
					hci_transport_h4_ecos.c \
					hci_transport_h5.c \
					l2cap.c \
					l2cap_signaling.c \
					classic/avdtp_acceptor.c \
					classic/avdtp_initiator.c \
					classic/avdtp_sink.c \
					classic/avdtp_source.c \
					classic/avdtp_util.c \
					classic/bnep.c \
					classic/btstack_cvsd_plc.c \
					classic/btstack_link_key_db_memory.c \
					classic/btstack_link_key_db_memory_save.c \
					classic/btstack_sbc_plc.c \
					classic/device_id_server.c \
					classic/hfp.c \
					classic/hfp_ag.c \
					classic/hfp_gsm_model.c \
					classic/hfp_hf.c \
					classic/hfp_msbc.c \
					classic/hsp_ag.c \
					classic/hsp_hs.c \
					classic/pan.c \
					classic/rfcomm.c \
					classic/sdp_client.c \
					classic/sdp_client_rfcomm.c \
					classic/sdp_server.c \
					classic/sdp_util.c \
					classic/spp_server.c \
					deamon/deamon.c \
					deamon/deamon_io.c 
                    
                    
    cdl_component CYGPKG_BLUETOOTH_CONFIG {
    	display		"Bluetooth library configuration."
    	flavor		none
    	description "
    		This component contans configuration option related to the
    		bluetooth stack."
    		
    	cdl_component CYGOPT_BLUETOOTH_ENABLE_BLE {
    		display 		"Enable support for BLE"
    		flavor			bool
    		default_value 	0
    		description "
    			This options enabes the bluetooth low energy
    			support in bluetooth stackt. NOTE: supoort for the
    			bluetooth low energy is not yet implmemented in
    			ecos bluetooth deamon."
    	}
    	
    	cdl_component CYGOPT_BLUETOOTH_ENABLE_CLASIC {
    		display 		"Enable support for classic bluetooth"
    		flavor			bool
    		default_value 	1
    		description "
    			This options enabes the clasic bluetooth
    			support in bluetooth stack."
    	}

    	cdl_component CYGPKG_BLUETOOTH_CONFIG_CLASIC {
    		display		"Configuratin for clasic bluetooth."
    		active_if    CYGOPT_BLUETOOTH_ENABLE_CLASIC
    		flavor		none
    	
	    	cdl_component CYGINT_BLUETOOTH_BNEP_SERVICES {
	    		display 		"Maximum BNEP services"
	    		active_if    CYGOPT_BLUETOOTH_ENABLE_CLASIC
	    		flavor			data
	    		default_value 	1
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum BNEP
	    			(Bluetooth Network Emulation Protocol) services."
	    	}
	    	
	    	cdl_component CYGINT_BLUETOOTH_HFP_CONNECTION {
	    		display 		"Maximum HFP connection"
	    		active_if    CYGOPT_BLUETOOTH_ENABLE_CLASIC
	    		flavor			data
	    		default_value 	0
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum HFP
	    			( Hands-Free Profile and Headset Profile) connections."
	    	}
	    	
	    	cdl_component CYGINT_BLUETOOTH_L2CAP_SERVICES {
	    		display 		"Maximum L2CAP services"
	    		active_if    CYGOPT_BLUETOOTH_ENABLE_CLASIC
	    		flavor			data
	    		default_value 	2
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum L2CAP services."
	    	}
	    	
	    	cdl_component CYGINT_BLUETOOTH_RFCOMM_SERVICES {
	    		display 		"Maximum RFCOMM services"
	    		active_if    CYGOPT_BLUETOOTH_ENABLE_CLASIC
	    		flavor			data
	    		default_value 	1
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum RFCOMM services."
	    	}
	    	
	    	cdl_component CYGINT_BLUETOOTH_SERVICE_RECORD_ITEMS {
	    		display 		"Maximum service records"
	    		active_if    CYGOPT_BLUETOOTH_ENABLE_CLASIC
	    		flavor			data
	    		default_value 	1
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum service records."
	    	}
	    	
	    	cdl_component CYGINT_BLUETOOTH_SPP_CONNECTIONS {
	    		display 		"Maximum SPP connections"
	    		active_if    CYGOPT_BLUETOOTH_ENABLE_CLASIC
	    		flavor			data
	    		default_value 	2
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum SPP(Serial Port Profile)
	    			entries."
	    	}
	    }
    	
    	cdl_component CYGPKG_BLUETOOTH_CONIG_BLE {
    		display		"Configuratin for ble bluetooth."
    		active_if    CYGOPT_BLUETOOTH_ENABLE_BLE
    		flavor		none
    		
	    	cdl_component CYGINT_BLUETOOTH_GATT_CLIENTS {
	    		display 		"Maximum GAT clients"
	    		active_if       CYGOPT_BLUETOOTH_ENABLE_BLE
	    		flavor			data
	    		default_value 	0
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum GATT
	    			(Generic Attribute Profile) clients."
	    	}
	    	
	    	cdl_component CYGINT_BLUETOOTH_GATT_SUB_CLIENTS {
	    		display 		"Maximum GAT sub-clients"
	    		active_if       CYGOPT_BLUETOOTH_ENABLE_BLE
	    		flavor			data
	    		default_value 	0
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum GATT
	    			(Generic Attribute Profile) sub-clients."
	    	}
	
	    	cdl_component CYGINT_BLUETOOTH_SM_LOOKUP_ENTRIES {
	    		display 		"Maximum sm lookup entris"
	    		active_if       CYGOPT_BLUETOOTH_ENABLE_BLE
	    		flavor			data
	    		default_value 	3
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum sm lookup entries."
	    	}
	    	
	    	cdl_component CYGINT_BLUETOOTH_WHITELIST_ENTRIES {
	    		display 		"Maximum whitelist entris"
	    		active_if       CYGOPT_BLUETOOTH_ENABLE_BLE
	    		flavor			data
	    		default_value 	1
	    		legal_values    0 to 10
	    		description "
	    			This options set maximum whitelist entries."
	    	}
    	}
    	
    	cdl_component CYGINT_BLUETOOTH_ACL_PAYLOAD_SIZE {
    		display 		"Maximum payload size "
    		flavor			data
    		default_value 	52
    		legal_values    52 to 2048
    		description "
    			This options set payload buffer size."
    	}
    	
    	cdl_component CYGPKG_BLUETOOTH_DEBUG_CONIG {
	    	display		"Bluetooth stack debug output configuration."
	    	flavor		none
	    	description " "
	    	
	    	cdl_component CYGOPT_BLUETOOTH_LOG_ERROR {
	    		display 		"Enable error output"
	    		flavor			bool
	    		default_value 	1
	    		description "
	    			This options enabes the to display error logs
	    			from the bluetooth stack."
	    	}
	    	
	    	cdl_component CYGOPT_BLUETOOTH_LOG_INFO {
	    		display 		"Enable info output"
	    		flavor			bool
	    		default_value 	1
	    		description "
	    			This options enabes the to display info logs
	    			from the bluetooth stack."
	    	}
	    	
	    	cdl_component CYGOPT_BLUETOOTH_LOG_DEBUG {
	    		display 		"Enable debug output"
	    		flavor			bool
	    		default_value 	0
	    		description "
	    			This options enabes the to display debug logs
	    			from the bluetooth stack."
	    	}
	    }
    }
    
    cdl_component CYGPKG_BLUETOOTH_DEAMON_CONIG {
    	display		"Bluetooth stack deamon configuration."
    	flavor		none
    	description " "
    	
    	cdl_component CYGOPT_BLUETOOTH_ECOS_DEAMON_ENABLE {
	    		display 		"Enable ecos bluetooth stack deamon."
	    		flavor			bool
	    		default_value 	1
	    		description "
	    			Enable ecos bluetooth stack deamon. Without ecos deamon
	    			it is possible to run native bleutooth stack applications."
	    }
	    
	    cdl_component CYGOPT_BLUETOOTH_ECOS_DEAMON_USE_RAD_QUEUE {
	    		display 		"Enable buffer for read oparation."
	    		active_if 		CYGOPT_BLUETOOTH_ECOS_DEAMON_ENABLE
	    		flavor			bool
	    		default_value 	1
	    		description "
	    			If this option is diabled it is not possible to receive data
	    			if something is porcessed."
	    }
	    
	    cdl_component CYGINT_BLUETOOTH_ECOS_DEAMON_RAD_QUEUE_SIZE {
	    		display 		"Size of the rad queue."
	    		active_if 		CYGOPT_BLUETOOTH_ECOS_DEAMON_ENABLE && CYGOPT_BLUETOOTH_ECOS_DEAMON_USE_RAD_QUEUE
	    		flavor			data
	    		default_value 	1024
	    		legal_values    64 to 65535
	    		description "
	    			Size of the read queue in bytes."
	    }
	    
	    cdl_component CYGINT_BLUETOOTH_ECOS_DEAMON_CHANNELS_COUNT {
	    		display 		"Number of the independednt bluetooth channels."
	    		active_if 		CYGOPT_BLUETOOTH_ECOS_DEAMON_ENABLE
	    		flavor			data
	    		default_value 	2
	    		legal_values    1 to 4
	    		description "
	    			This options depends as well on bluetooths stack channel configurations.
	    			For naw only 4 channels can be used."
	    }
	    
	    cdl_component CYGINT_BLUETOOTH_ECOS_DEAMON_STORE_LINK_KEY_TO_MEMORY {
	    		display 		"Store link keys to ram storage."
	    		active_if 		CYGOPT_BLUETOOTH_ECOS_DEAMON_ENABLE
	    		flavor			bool	
	    		default_value 	1
	    		description "
	    			If htis option is enabled the link keys asre store to
	    			ram storage. If this option is disabled the keys are
	    			stored to permanent memory. Permanent storage is not 
	    			yet universally implemented."
	    }
	    
	    cdl_component CYGINT_BLUETOOTH_ECOS_DEAMON_LOCAL_NAME {
	    		display 		"Name of the bluetooth device."
	    		active_if 		CYGOPT_BLUETOOTH_ECOS_DEAMON_ENABLE
	    		flavor			data	
	    		default_value 	{"\"eCos\""}
	    		description "
	    			If htis option sets the name of the bluetooth device."
	    }
	    
    }
}

# ====================================================================
# End of bluetooth.cdl
