# ====================================================================
#
#      lua.cdl
#
#      Lua
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Mike Jones <mike@proclivis.com>
# Contributors:
# Date:           2014-01-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_LUA {
    display       "Lua language support"
    description   "
            This component supports running Lua scripts."
    doc           doc/manual.html
    include_dir   cyg/lua
    requires      CYGPKG_ISOINFRA
    compile       lapi.c lcode.c ldebug.c lgc.c lmathlib.c lopcodes.c 
    compile       lstring.c ltm.c lvm.c lauxlib.c lcorolib.c ldo.c linit.c 
    compile       lmem.c loslib.c lstrlib.c lua.c lzio.c lbaselib.c lctype.c
    compile       ldump.c liolib.c loadlib.c lparser.c ltable.c luac.c lbitlib.c
    compile       ldblib.c lfunc.c llex.c lobject.c lstate.c ltablib.c lundump.c

# ====================================================================

    cdl_option CYGPKG_LUA_CFLAGS_ADD {
        display "Additional compiler flags"
        flavor  data
        no_define
        default_value { "-DLUA_USE_POSIX" }
        description   "
	    This option modifies the set of compiler flags for
	    building this package. These flags are used in addition
	    to the set of global flags."
    }
    
    cdl_option CYGPKG_LUA_ROOT {
        display "Root directory"
        flavor  data
        default_value { "\"/disk0/usr/local/\"" }
        description   "
	    This option sets the root direcotry of the file system 
	    and the base directory for lua files."
    }

}

# ====================================================================
# EOF lua.cdl
