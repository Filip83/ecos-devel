##==========================================================================
##
##      adc_ltc2498_freescale_dspi.cdl
##
##      LTC2498 ADC instatntiation for Freescale DSPI
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                  
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Mike Jones
## Date:         2013-06-12
##
######DESCRIPTIONEND####
##
##==========================================================================

cdl_package CYGPKG_DEVS_ADC_LTC2498_FREESCALE_DSPI {
    display "Driver for LTC2498 adc over Freescale DSPI"
    parent CYGPKG_DEVS_ADC_SPI_LTC2498
    
    cdl_component CYGHWR_DEVS_ADC_SPI_LTC2498_DEV0 {
        display "Use LTC2498 ADC device 0"
        flavor bool
        default_value 0
        no_define
        
        requires CYGPKG_DEVS_ADC_SPI_LTC2498
        requires CYGPKG_DEVS_SPI_FREESCALE_DSPI
        implements CYGHWR_DEVS_ADC_SPI_LTC2498_DEVICE
        
        requires CYGHWR_DEVS_ADC_LTC2498_DEV0_SPI_BUS
        requires CYGHWR_DEVS_ADC_LTC2498_DEV0_SPI_CS == 1
        
        compile -library=libextras.a adc_ltc2498_freescale_dspi.c
        
        cdl_component CYGHWR_DEVS_ADC_LTC2498_DEV0_SPEED {
            display "Nominal clock speed Hz"
            flavor data
            default_value 2000000
            
            cdl_option CYGHWR_DEVS_ADC_LTC2498_DEV0_SPI_USE_DBR {
                display "Use double baud rate"
                flavor bool
                default_value 0
                description "
                    Double baud rate is a feature of Freescale DSPI
                    that may provide higher baud rates but duty the cycle may be
                    different than 50/50 depdent on scaler/prescaler setting
                    for achieved baud rate."
            }
        }
        
        cdl_option CYGHWR_DEVS_ADC_LTC2498_DEV0_CS_DLY {
            display "Nominal chip select delays (units)"
            flavor data
            legal_values { 1 10 }
            default_value 1
        }
        
        cdl_option CYGHWR_DEVS_ADC_LTC2498_DEV0_CS_DLY_UN {
            display "Chip select delay unit (ns)"
            flavor data
            default_value 100
            legal_values { 100 1000 }
        }
    }
}
