# ====================================================================
#
#      hal_avr32_km_8.cdl
#
#      AVR32 Platform HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Original data:  
# Contributors:
# Date:           2016-05-09
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_AVR32_KM_8 {
    display  "KM-8 board"
    parent        CYGPKG_HAL_AVR32
    include_dir   cyg/hal
    hardware
    description   "
           The AVR32 HAL package should be used when targetting the
           AVR32 Platform."

    compile       hal_diag.c hal_aux.c gpio.c board_config.c pcf_wallclock.c

    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_avr32.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_avr32_km_8.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_BOARD_H    <cyg/hal/board_config.h>"
        puts $::cdl_system_header "#define CYGHWR_MEMORY_LAYOUT_H <pkgconf/mlt_avr32_uc3c.h>"
        puts $::cdl_system_header "#define CYGHWR_MEMORY_LAYOUT_LDI <pkgconf/mlt_avr32_uc3c.ldi>"
    }

     cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor none
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator(Not realy used)"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value {CYGHWR_HAL_AVR32_CPU_FREQ * 1000000 / CYGNUM_HAL_RTC_DENOMINATOR}
            description   "
                The tick timer facility is used
                to drive the eCos kernel RTC. The count register
                increments at the CPU clock speed.  By default, 100 Hz"
        }
    }

   # CPU clk specifics
    cdl_component CYGNUM_HAL_CLOCK_CONSTANTS {
        display       "CPU clock constants."
        flavor        none

        cdl_option CYGNUM_HAL_MAIN_CLOCK_SOURCE {
            display       "Select main clock source"
            flavor        data
            legal_values  { "RCSYS" "OSC0" "DFLL" "RC120M" }
            default_value { "RC120M"}
        }
        cdl_option CYGNUM_HAL_CPU_CLOCK_DIVIDER {
            display       "CPU clock divider 2^(value + 1)"
            flavor        booldata
            legal_values  0 to 8
            default_value 0
        }

	cdl_option CYGNUM_HAL_PBA_CLOCK_DIVIDER {
            display       "PBA domain clock divider 2^(value + 1)"
            flavor        booldata
            legal_values  0 to 8
            default_value 0
        }

	cdl_option CYGNUM_HAL_PBB_CLOCK_DIVIDER {
            display       "PBB domain clock divider 2^(value + 1)"
            flavor        booldata
            legal_values  0 to 8
            default_value 0
        }
    }

    # CPU oscilators specifics
    cdl_component CYGNUM_HAL_OSCILATORS_CONSTANTS {
        display       "Oscilators constants."
        flavor        none

	cdl_component CYGNUM_HAL_OSCILATORS_OSC0_CONSTRAINS {
            display       "Oscilator 0 settings"
            flavor        none
            
		cdl_option CYGNUM_HAL_OSCILATORS_OSC0_ENABLED {
		    display       "Enable osciloator 0"
		    flavor        bool
		    default_value 1
		}
		
		cdl_option CYGNUM_HAL_OSCILATORS_OSC0_FREQV {
		    display       "Osciloator 0 frequency MHz"
		    flavor        data
		    default_value 16
		    active_if  CYGNUM_HAL_OSCILATORS_OSC0_ENABLED
		}


		cdl_option CYGNUM_HAL_OSCILATORS_OSC0_AGC_ENABLE {
		    display       "Osciloator 0 AGC enable"
		    flavor        bool
		    default_value 1
		    active_if  CYGNUM_HAL_OSCILATORS_OSC0_ENABLED
		}

		cdl_option CYGNUM_HAL_OSCILATORS_OSC0_CRYSTAL {
		    display       "Osciloator 0 crystal."
		    flavor        bool
		    default_value 1
		    active_if  CYGNUM_HAL_OSCILATORS_OSC0_ENABLED
		}

		cdl_option CYGNUM_HAL_OSCILATORS_OSC0_EXTERNAL_STARTUP_TIME {
		    display       "Osciloator 0 external source startup time"
		    flavor        data
		    legal_values  0 to 14
		    default_value 14
		    active_if CYGNUM_HAL_OSCILATORS_OSC0_EXTERNAL
		}
            }

            #-------------
            cdl_component CYGNUM_HAL_OSCILATORS_OSC32K_CONSTRAINS {
                display       "32kHz oscilator settings"
                flavor        none

                    cdl_option CYGNUM_HAL_OSCILATORS_OSC32K_ENABLED {
                        display       "Enable 32kHz osciloator"
                        flavor        bool
                        default_value 1
                    }

                    cdl_option CYGNUM_HAL_OSCILATORS_OSC32K_EXTERNAL {
                        display       "32kHz oscilator use external source"
                        flavor        bool
                        default_value 0
                        active_if  CYGNUM_HAL_OSCILATORS_OSC32K_ENABLED
                    }

                    cdl_option CYGNUM_HAL_OSCILATORS_OSC32K_MODE {
                        display       "32kHz oscilator normal I-current mode"
                        flavor        bool
                        default_value 1
                        active_if  !CYGNUM_HAL_OSCILATORS_OSC32K_EXTERNAL
                    }

                    cdl_option CYGNUM_HAL_OSCILATORS_OSC32K_EXTERNAL_STARTUP_TIME {
                        display       "Osciloator 1 external source startup time"
                        flavor        data
                        legal_values  0 to 7
                        default_value 4
                        active_if CYGNUM_HAL_OSCILATORS_OSC32K_EXTERNAL
                    }
                }		

                #-------------
                cdl_component CYGNUM_HAL_OSCILATORS_RC120M_CONSTRAINS {
                    display       "120MHz oscilator settings"
                    flavor        none

                        cdl_option CYGNUM_HAL_OSCILATORS_RC120M_ENABLED {
                            display       "Enable 120MHz internal rc osciloator"
                            flavor        bool
                            default_value 1
                        }
                }	

                #-------------
                cdl_component CYGNUM_HAL_OSCILATORS_RC32K_CONSTRAINS {
                    display       "32kHz internal RC oscilator settings"
                    flavor        none

                        cdl_option CYGNUM_HAL_OSCILATORS_RC32K_ENABLED {
                            display       "Enable 32kHz internal rc osciloator"
                            flavor        bool
                            default_value 0
                        }
                }	

	#-------------
	cdl_component CYGNUM_HAL_OSCILATORS_PLL0_CONSTRAINS {
            display       "PLL0 settings"
            flavor        none
            
		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_ENABLED {
		    display       "Enable PLL0"
		    flavor        bool
		    default_value 1
		}

		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_SOURCE {
		    display       "Select PLL0 clock source"
		    flavor        data
		    legal_values  { "OSC0" "GCLK8"}
		    default_value { "OSC0"}
		}
		
		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_DIVIDER {
		    display       "PLL0 divider"
		    flavor        data
		    legal_values 0 to 15
		    default_value 2
		}
		
		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_MULTIPLIER {
		    display       "PLL0 multiplier"
		    flavor        data
		    legal_values 0 to 15
		    default_value 5
		}

		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_START_COUNT {
		    display       "PLL start up time."
		    flavor        data
		    legal_values 0 to 63
		    default_value 10
                    description "Specifies the number of RCSYS clock cycles 
                    before ISR.PLLLOCKn will be set after PLLn has been written, 
                    or after PLLn has been automatically re-enabled after 
                    exiting a sleep mode."
		}

		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_VCO_FREQ {
		    display       "PLL0 VCO frequency range"
		    flavor        bool
		    default_value 0
		}
		
		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_OUTPUT_DIVIDER {
		    display       "Enable additional output divder (2)"
		    flavor        bool
		    default_value 0
		}

		cdl_option CYGNUM_HAL_OSCILATORS_PLL0_BANDWIDTH_MODE {
		    display       "Dsable wide bandwidth mode"
		    flavor        bool
		    default_value 0
		}
	}


	#-------------
	cdl_component CYGNUM_HAL_OSCILATORS_DFLL0_CONSTRAINS {
            display       "DFLL0 settings"
            flavor        none
            
		cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_ENABLED {
		    display       "Enable DFLL0"
		    flavor        bool
		    default_value 0
		}

                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_MODE {
		    display       "Select open loop or cloded loop operation."
		    flavor        bool
		    default_value 1
                    description "If this option is enabled closed llop mode is
                                selected, open loop mode otherwise"
		}

                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_DITHERING {
		    display       "Enable dithering mode."
		    flavor        bool
		    default_value 1
                    active_if      CYGNUM_HAL_OSCILATORS_DFLL0_MODE == 1
		}
                
                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_LLAW {
		    display       "Enable lose of clock after wakeup."
		    flavor        bool
		    default_value 0
		}

                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_CCEN {
		    display       "Enable chill cycle."
		    flavor        bool
		    default_value 0
		}
                
                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_QLEN {
		    display       "Enable quick lock."
		    flavor        bool
		    default_value 1
                    active_if      CYGNUM_HAL_OSCILATORS_DFLL0_MODE == 1
		}

                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_FINE_MAX_STEPP {
		    display       "FINE Calibration Value"
		    flavor        data
		    legal_values  0 to 511
		    default_value 4
                    active_if      CYGNUM_HAL_OSCILATORS_DFLL0_MODE == 1
		}
                
                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_COARSE_MAX_STEPP {
		    display       "Coarse Calibration Value"
		    flavor        data
		    legal_values  0 to 255
		    default_value 4
                    active_if      CYGNUM_HAL_OSCILATORS_DFLL0_MODE == 1
		}

		cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_SOURCE {
		    display       "Select PLL1 clock source"
		    flavor        data
		    legal_values  { "RCSYS" "OSC32K" "OSC0"
                                    "RS120M" "CLKCPU" "RC32K" 
                                    "CLK1K"
                                  }
		    default_value { "OSC0"}
		}
		
                cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_DITHERING_SOURCE {
		    display       "Select dithering clock source"
		    flavor        data
		    legal_values  { "RCSYS" "OSC32K" "OSC0"
                                    "RS120M" "CLKCPU" "RC32K" 
                                    "CLK1K"
                                    "PLL0" "GCLKIN0" "GCLKIN1"
                                    "GCLKIN2" "GCLK9"
                                  }
		    default_value { "OSC0"}
                    active_if      CYGNUM_HAL_OSCILATORS_DFLL0_DITHERING == 1
		}
		

		cdl_option CYGNUM_HAL_OSCILATORS_DFLL0_FREQ {
		    display       "DFLL output frequency in kHz"
                    flavor  data
		    legal_values 0.0001 to 50000.0000
                    default_value 23961.6
		}
	}
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        description   "
            Global build options including control over
            compiler flags, linker flags and choice of toolchain."


        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "avr32" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS .
                            "-mpart=uc256l3u -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions "
            }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-mpart=uc256l3u -Wl,--gc-sections -Wl,-static -g -nostdlib"  }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_option CYGHWR_HAL_AVR32_CPU_FREQ {
        display "CPU frequency"
        flavor  data
        legal_values 0.0001 to 50.0000
        default_value 23.9616
        description "
           This option contains the frequency of the CPU in MegaHertz.
           Choose the frequency to match the processor you have. This
           may affect thing like serial device, interval clock and
           memory access speed settings."
    }

    cdl_option CYGHWR_RAM_SIZE {
        display       "Size of RAM memory"
        flavor        data
        default_value 0x10000
        description   "
            Size of RAM memory. This value is used to generate linker script.
            Not used yet."
    }

    cdl_option CYGHWR_ROM_SIZE {
        display       "Size of ROM memory"
        flavor        data
        default_value 0x80000
        description   "
            Size of ROM memory. This value is used to generate linker script.
            Not used yet."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200 230400
        default_value 57600
        description   "
            This option selects the baud rate used for the diagnostic console.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same.
            Note: very high baud rates are useful during simulation."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200 230400
        default_value 57600
        description   "
            This option controls the baud rate used for the GDB connection.
            Note: very high baud rates are useful during simulation."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        default_value  5
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The ORP platform has at least one serial port, but it can potentially have several.
           This option chooses which port will be used to connect to a host
           running GDB."
    }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    2
        description      "
           The ORP platform has at least one serial port, but it can potentially have several.
           This option chooses which port will be used for diagnostic output."
     }

    define_proc {
        puts $cdl_header "#define CYGHWR_HAL_VSR_TABLE    0"
        puts $cdl_header "#define CYGHWR_HAL_VIRTUAL_VECTOR_TABLE 0xF00"
    }
}

# EOF hal_avr32_km_8.cdl
