##==========================================================================
##
##      kinetis_clocking.cdl
##
##      Cortex-M Freescale Kinetis Clocking
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Ilija Kocho <ilijak@siva.com.mk>
## Date:         2011-10-19
##
######DESCRIPTIONEND####
##
##==========================================================================


#    cdl_component CYGHWR_HAL_CORTEXM_KINETIS_CLOCKING
#    display       "Clocking"

    cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ {
        display "System frequency actual value"
        flavor data
        calculated { CYGNUM_HAL_CORTEXM_KINETIS_MCG_MCGOUT_FREQ_SP  }
        description "Operating system clock frequency."
    }

    cdl_component CYGHWR_HAL_CORTEXM_KINETIS_MCG {
        display "MCG"
        flavor data
        no_define
        calculated { CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK . " " .
            ((CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ+500000)/1000000) . "MHz, " . (
                  (CYGOPT_HAL_CORTEXM_KINETIS_MCG_FLL_PLL_REFSRC == "EXT_REFCLK") ?
                  CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS :
                  CYGOPT_HAL_CORTEXM_KINETIS_MCG_FLL_PLL_REFSRC)

        }
        description "Multipurpose Clock Generator"

        cdl_option CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK {
            display "System clock source"
            flavor data
            default_value { "FLL" }
            legal_values {
                "PLL" "FLL" "EXT_REFCLK" "INT_RC"
            }
            requires { CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "PLL" implies
                CYGOPT_HAL_CORTEXM_KINETIS_MCGOUT_PLL == 1
            }
            description "
                Select one of 4 options for MCG output clock:
                PLL, FLL oscillator, External reference clock or internal
                RC oscilator."
        }

        cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_MCGOUT_FREQ_SP {
                display "MCGOUT output frequency set point"
                flavor data
                legal_values  32768 to 1200000000
                calculated {
                    (CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "FLL") ? 
                       CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_FREQ_AV :
                    (CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "PLL") ? 
                     CYGNUM_HAL_CORTEXM_KINETIS_100_MCG_PLL_FREQ_AV :
                    (CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "EXT_REFCLK") ?
                     CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ :
                     CYGOPT_HAL_CORTEXM_KINETIS_MCGOUT_INT_RC
                }
                description "MCGOUT output frequency."

        }

        cdl_component CYGOPT_HAL_CORTEXM_KINETIS_MCG_OSC0 {
            display "OSC0 source clock settings"
            flavor bool
            default_value 1
            description "Configure OSC0 paramters."

            cdl_option CYGOPT_HAL_CORTEXM_KINETIS_MCG_OSC0_IS {
                display "Clock type"
                flavor data
                default_value { "OSC" }
                legal_values { "OSC" "XTAL" }

                requires {
                    (CYGOPT_HAL_CORTEXM_KINETIS_MCG_OSC0_IS == "OSC") implies
                    (CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ <= 50000000)
                }

                requires {
                    (CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL") implies
                    (((CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ >= 3000000) &&
                      (CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ <= 32000000)) ||
                      ((CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ >= 32000) &&
                       (CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ <= 40000)))
                }

                description "
                Ext reference can be External oscillator or a crystal
                for the on-chip oscillator."
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ {
                display "Clock frequency"
                flavor data
                legal_values  0 to 50000000
                default_value 4000000
                description "External oscillator or crystal reference in Hz."
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_OSC_CAP {
                display "XTAL parallel C \[pF\]"
                flavor data
                active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_REF_EXT_IS == "XTAL" }
                legal_values { 0 2 4 6 8 10 12 14 16 18 20 22 24 26 28 30 32 }
                default_value { 0 }
                description "
                    The oscillator has 4 on-chip capacitors that combined
                    produce capacitance in parallel to the crystal."
                }
        }

        cdl_component CYGOPT_HAL_CORTEXM_KINETIS_MCGOUT_FLL {
            display "FLL oscillator"
            flavor none
            no_define
            active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "FLL" }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_SOURCE {
                display "Reference frequency source"
                flavor data
                legal_values { "INTERNAL_32K" "EXT_OSC0" "EXT_32K_RTC" "EXT_OSC1" }
                default_value { "INTERNAL_32K" }

                requires {
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_SOURCE == "EXT_OSC0") implies
                      CYGOPT_HAL_CORTEXM_KINETIS_MCG_OSC0 == 1 
                         }

            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_REF_FREQ {
                display "DCO input frequency"
                flavor data
                calculated {
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_SOURCE == "INTERNAL_32K" ||
                     CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_SOURCE == "EXT_32K_RTC") ?
                    32765 :  CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ
                }
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_RANGE {
                display "Reference frequency range"
                flavor data
                legal_values 0 1 2
                default_value { 
                (CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_SOURCE == "INTERNAL_32K" ||
                 CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_SOURCE == "EXT_32K_RTC") ? 0 :
                (CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_SOURCE == "EXT_OSC0") ?
                 ((CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_REF_FREQ >= 40000) ? 1 : 0) : 1 
                             }          
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FRDIV_REG {
                display "FLL divider register value"
                flavor data
                legal_values 0 1 2 3 4 5 6 7
                default_value 0
            }

            cdl_option CYGNUM_HAL_CORTEXM_MCG_DCO_DRST_DRS {
                display "DCO Range Select"
                flavor data
                legal_values 0 1 2 3
                default_value {
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_PLL_FREQ_SP) >= 80000000 ? 3 :
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_PLL_FREQ_SP) >= 60000000 ? 2 :
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_PLL_FREQ_SP) >= 40000000 ? 1 : 0
                }
            }

            cdl_option CYGNUM_HAL_CORTEXM_MCG_DCO_DMX32 {
                display "DCO max. frequency with 32768 reference"
                flavor data
                legal_values { 0 0x80 }
                default_value { 0x80}
            }

            cdl_option CYGNUM_HAL_CORTEXM_MCG_DCO_FLL_FACT {
                display "FLL factor"
                flavor data
                calculated {
                    (CYGNUM_HAL_CORTEXM_MCG_DCO_DMX32 == 0x80) ?
                    ((CYGNUM_HAL_CORTEXM_MCG_DCO_DRST_DRS == 0 ) ?  732 :
                     (CYGNUM_HAL_CORTEXM_MCG_DCO_DRST_DRS == 1 ) ? 1464 :
                     (CYGNUM_HAL_CORTEXM_MCG_DCO_DRST_DRS == 2 ) ? 2197 : 2929 ) :
                    ((CYGNUM_HAL_CORTEXM_MCG_DCO_DRST_DRS == 0 ) ?  640 :
                     (CYGNUM_HAL_CORTEXM_MCG_DCO_DRST_DRS == 1 ) ? 1280 :
                     (CYGNUM_HAL_CORTEXM_MCG_DCO_DRST_DRS == 2 ) ? 1920 : 2560 )
                }
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_DCO_IN {
                display "DCO input frequency"
                flavor data
                calculated { CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_REF_FREQ /
                    ( CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FRDIV_REG == 0 ?
                     ((CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_RANGE == 0) ? 1 : 32 ) :
                     (CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FRDIV_REG *
                      ((CYGNUM_HAL_CORTEXM_KINETIS_MCG_REF_FREQ_RANGE == 0) ? 2 : 64)))
                }
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_DCO_IN_CHECK {
                display "DCO input frequency check"
                flavor data
                no_define
                legal_values { "OK" "NOK" "not applicable" }
                calculated {
                    CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "FLL" ?
                    ((CYGNUM_HAL_CORTEXM_KINETIS_MCG_DCO_IN >= 31250) &&
                     (CYGNUM_HAL_CORTEXM_KINETIS_MCG_DCO_IN <= 39063) ?
                     "OK" : "NOK" ) :
                    "NotApplicable"
                }
                active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "FLL" }
                requires {
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_DCO_IN >= 31250) &&
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_DCO_IN <= 39063)
                }
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_FLL_FREQ_AV {
                display "FLL output frequency actual value"
                flavor data
                calculated {CYGNUM_HAL_CORTEXM_KINETIS_MCG_DCO_IN *
                    CYGNUM_HAL_CORTEXM_MCG_DCO_FLL_FACT }
            }
        }

        cdl_component CYGOPT_HAL_CORTEXM_KINETIS_MCGOUT_PLL {
            display "PLL oscillator"
            flavor none
            no_define
            active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK == "PLL" &&
                        CYGOPT_HAL_CORTEXM_KINETIS_MCG_OSC0 == 1 }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ {
                display "PLL input frequency"
                flavor data
                calculated { CYGHWR_HAL_CORTEXM_KINETIS_MCG_OSC0_FREQ }
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_INFREQ_X {
                display "Phase detector proposed input frequency"
                no_define
                flavor data
                calculated {
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ > 180000000) ?
                    3800000 :
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ > 110000000) ?
                    3000000 :
                    !(CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ % 3) ? 2000000 :
                    !(CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ % 4) ? 2000000 :
                    !(CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ % 5) ? 2500000 :
                    300000
                }
            }

            cdl_option CYGOPT_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_PRDIV {
                display "PLL External Reference Divider"
                flavor data
                legal_values 1 to 24
                default_value {
                    CYGNUM_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_INFREQ_X ?
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ /
                     CYGNUM_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_INFREQ_X ) : -1
                }
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_INFREQ {
                display "Phase detector input frequency"
                no_define
                flavor data
                legal_values 2000000 to 4000000
                calculated { CYGOPT_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_PRDIV ?
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ /
                     CYGOPT_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_PRDIV) : -1
                }
            }

            cdl_option CYGOPT_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_VDIV {
                display "VCO Divider"
                flavor data
                legal_values 24 to 55
                default_value 24
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_100_MCG_PLL_FREQ_AV {
                display "PLL output frequency actual value"
                flavor data
                calculated { CYGOPT_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_PRDIV ?
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCG_PLL_REF_FREQ /
                     CYGOPT_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_PRDIV *
                     CYGOPT_HAL_CORTEXM_KINETIS_100_MCGOUT_PLL_VDIV) : -1
                }
            }
        }
        

        cdl_component CYGOPT_HAL_CORTEXM_KINETIS_MCGOUT_INT_RC {
            display "Internal Reference Clock"
            flavor data
            calculated { CYGOPT_HAL_CORTEXM_KINETIS_MCGOUT_INT_RC_HI ? 4000000 : 32768 }
            active_if { CYGOPT_HAL_CORTEXM_KINETIS_MCG_MCGOUTCLK ==  "INT_RC" }

            cdl_option CYGOPT_HAL_CORTEXM_KINETIS_MCGOUT_INT_RC_HI {
                display "Use highh frequency internal osc."
                flavor bool
                default_value 1
            }
        }
    }

    cdl_component CYGHWR_HAL_CORTEXM_KINETIS_CLK_DIST {
        display "Subsystem clocking"
        flavor none
        no_define

        cdl_component CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_BUS {
            display "Peripheral bus"
            flavor data
            calculated { CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                CYGHWR_HAL_CORTEXM_KINETIS_CLKDIV_PER_BUS
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_MAX {
                display "Frequency limit"
                flavor data
                default_value 50000000
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_BUS_SP {
                display "Calculated value"
                flavor data
                default_value {
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ <=
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_MAX ?
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ :
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_MAX
                }
                legal_values  0 to CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_MAX
            }
            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLKDIV_PER_BUS {
                display "Divider"
                flavor data
                legal_values 1 to 16

                default_value { !(CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ %
                                  CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_BUS_SP)  ?
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                     CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_BUS_SP)  :
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                     CYGHWR_HAL_CORTEXM_KINETIS_CLK_PER_BUS_SP + 1)
                }
            }
        }

        cdl_component CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH {
            display "Flash"
            flavor data
            calculated { CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                CYGHWR_HAL_CORTEXM_KINETIS_CLKDIV_FLASH
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_MAX {
                display "Frequency limit"
                flavor data
                default_value 25000000
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_SP {
                display "Calculated value"
                flavor data
                default_value {
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ <=
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_MAX ?
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ :
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_MAX
                }
                legal_values  0 to CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_MAX
            }
            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLKDIV_FLASH {
                display "Divider"
                flavor data
                legal_values 1 to 16

                default_value {
                    !(CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ %
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_SP)  ?
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                     CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_SP)  :
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                     CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLASH_SP + 1)
                }
            }
        }

        cdl_component CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS {
            display "Flex bus"
            flavor data
            calculated { CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                CYGHWR_HAL_CORTEXM_KINETIS_CLKDIV_FLEX_BUS
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_MAX {
                display "Frequency limit"
                flavor data
                default_value 50000000
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_SP {
                display "Calculated value"
                flavor data
                default_value {
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ <=
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_MAX ?
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ :
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_MAX
                }
                legal_values  0 to CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_MAX
            }
            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLKDIV_FLEX_BUS {
                display "Divider"
                flavor data
                legal_values 1 to 16

                default_value {
                    !(CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ %
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_SP)  ?
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                     CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_SP)  :
                    (CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ /
                     CYGHWR_HAL_CORTEXM_KINETIS_CLK_FLEX_BUS_SP + 1)
                }
            }
        }


        cdl_component CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB {
            display "USB clock"
            flavor data
            calculated { CYGNUM_HAL_CORTEXM_KINETIS_CLK_USB_IN *
                CYGHWR_HAL_CORTEXM_KINETIS_USBCLK_FRAC /
                CYGHWR_HAL_CORTEXM_KINETIS_USBCLK_DIV
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_MAX {
                display "Frequency limit"
                flavor data
                default_value 48000000
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_USBCLK_FRAC {
                display "Fractional Divider"
                flavor data
                legal_values 1 to 2
                default_value {
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ <
                    CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_MAX ? 1 :
                    ((CYGNUM_HAL_CORTEXM_KINETIS_CLK_USB_IN) >
                     (CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_SP * 4) ? 1 :
                     (CYGNUM_HAL_CORTEXM_KINETIS_CLK_USB_IN %
                      CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_SP ? 2 : 1))
                }
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_USBCLK_DIV {
                display "Divider"
                flavor data
                legal_values 1 to 8
                default_value { !((CYGNUM_HAL_CORTEXM_KINETIS_CLK_USB_IN *
                                   CYGHWR_HAL_CORTEXM_KINETIS_USBCLK_FRAC) %
                                   CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_SP)  ?
                    (CYGNUM_HAL_CORTEXM_KINETIS_CLK_USB_IN *
                     CYGHWR_HAL_CORTEXM_KINETIS_USBCLK_FRAC /
                     CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_SP)  :
                    ((CYGNUM_HAL_CORTEXM_KINETIS_CLK_USB_IN *
                      CYGHWR_HAL_CORTEXM_KINETIS_USBCLK_FRAC /
                      CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_SP) +1)
                }
            }

            cdl_option CYGNUM_HAL_CORTEXM_KINETIS_CLK_USB_IN {
                display "USB divider input frequency"
                flavor data
                calculated {
                    CYGNUM_HAL_CORTEXM_KINETIS_MCGOUT_FREQ
                }
            }

            cdl_option CYGHWR_HAL_CORTEXM_KINETIS_CLK_USB_SP {
                display "Desired"
                flavor data
                calculated 48000000
            }
        }

        cdl_option CYGHWR_HAL_CORTEXM_KINETIS_TRACECLK {
            display "Trace clock source"
            flavor data
            default_value { "CORE" }
            legal_values { "CORE" "MCGOUT" }

        }
        cdl_option CYGHWR_HAL_CORTEXM_KINETIS_TRACE_CLKOUT {
            display "Enable Trace Clock out"
            flavor bool
            default_value 0
        }
    }

    cdl_interface CYGINT_HAL_CORTEXM_KINETIS_RTC {
        display "System uses Real Time Clock"
    }

    cdl_component CYGHWR_HAL_CORTEXM_KINETIS_RTC {
        display "Real Time Clock"
        flavor bool
        default_value CYGINT_HAL_CORTEXM_KINETIS_RTC


        cdl_option CYGHWR_HAL_CORTEXM_KINETIS_RTC_OSC_CAP {
            display "RTC XTAL parallel C \[pF\]"
            flavor data
            legal_values { 0 2 4 6 8 10 12 14 16 18 20 22 24 26 28
                30 32 }
            default_value 0
            description "
                The Real Time Clock oscillator has 4 capacitors that
                combined produce capacitance in parallel to the crystal."
        }
    }

    # EOF kinetis_clocking.cdl
