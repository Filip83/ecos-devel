# ====================================================================
#
#      hal_arm_wandboard.cdl
#
#      Freescake i.MX6 Wandboard package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2006 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Mike Jones
# Contributors:
# Date:           2013-08-08
#
#####DESCRIPTIONEND####

cdl_package CYGPKG_HAL_ARM_IMX6_WANDBOARD {

    display       "Freescale Wandboard"
    parent         CYGPKG_HAL_ARM_IMX6

    include_dir    cyg/hal
    define_header  hal_arm_wandboard.h
    hardware

    description    "
        This HAL platform package provides generic
        support for the Freescale Wandboard."

    compile       wandboard_misc.c platform_init.c cortexA9.S

    implements    CYGINT_HAL_ARM_ARCH_ARM_CORTEXA9

    implements    CYGINT_IO_SERIAL_FREESCALE_UART0
    implements    CYGINT_HAL_FREESCALE_UART0
    implements    CYGINT_IO_FREESCALE_I2CA0
    implements    CYGINT_IO_FREESCALE_I2CA1
    implements    CYGINT_IO_FREESCALE_I2CA2

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_imx6.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_wandboard.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"Cortex-A9\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Freescale Wandboard\""
#        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { 
		(CYG_HAL_STARTUP == "RAM") ? 
			"arm_wandboard_ram" : 
			(CYG_HAL_STARTUP == "SD") ? 
				"arm_wandboard_sd" : 
				"arm_wandboard_rom" 
	    }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { 
		    (CYGPKG_HAL_SMP_CPU_MAX == 2) ?
			    ((CYGBLD_BUILD_REDBOOT) ? 
				    "<pkgconf/mlt_arm_wandboard_redboot_2.ldi>" : 
				    (CYG_HAL_STARTUP == "RAM") ? 
					    "<pkgconf/mlt_arm_wandboard_ram_2.ldi>" : 
					    "<pkgconf/mlt_arm_wandboard_sd_2.ldi>") :
		    ((CYGBLD_BUILD_REDBOOT) ? 
			    "<pkgconf/mlt_arm_wandboard_redboot_4.ldi>" : 
			    (CYG_HAL_STARTUP == "RAM") ? 
				    "<pkgconf/mlt_arm_wandboard_ram_4.ldi>" : 
				    "<pkgconf/mlt_arm_wandboard_sd_4.ldi>")
	        }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { 
		    (CYGPKG_HAL_SMP_CPU_MAX == 2) ?
			    ((CYGBLD_BUILD_REDBOOT) ? 
				    "<pkgconf/mlt_arm_wandboard_redboot_2.h>" : 
				    (CYG_HAL_STARTUP == "RAM") ? 
					    "<pkgconf/mlt_arm_wandboard_ram_2.h>" : 
					    "<pkgconf/mlt_arm_wandboard_sd_2.h>") :
		    ((CYGBLD_BUILD_REDBOOT) ? 
			    "<pkgconf/mlt_arm_wandboard_redboot_4.h>" : 
			    (CYG_HAL_STARTUP == "RAM") ? 
				    "<pkgconf/mlt_arm_wandboard_ram_4.h>" : 
				    "<pkgconf/mlt_arm_wandboard_sd_4.h>")
	        }
        }

	    cdl_option CYGHWR_MEMORY_LAYOUT_SD {
            display "Include SD Data in build"
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_SD
            flavor bool
            calculated { (CYG_HAL_STARTUP == "SD") }
        }
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display       "Number of communication channels on the board"
        flavor        data
        calculated    1
        description   "
            The wandboard SD has one serial port: UART0."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The wandboard SD has two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description      "
            The wandboard SD board has two UART serial ports. This option
            chooses which port will be used for diagnostic output."
     }
     
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        description   "
            This option selects the baud rate used for the diagnostic port."
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
         display       "GDB serial port baud rate"
         flavor        data
         legal_values  9600 19200 38400 57600 115200
         default_value 38400
         description   "
            This option controls the baud rate used for the GDB connection."
     }

    cdl_option CYGHWR_FREESCALE_ENET_MII_MDC_HAL_CLOCK {
        display "ENET MII MDC clock provided by HAL"
        flavor data
        active_if CYGPKG_DEVS_ETH_FREESCALE_ENET
        parent CYGPKG_DEVS_ETH_FREESCALE_ENET
        calculated 66000000
        description "
            ENET needs a clock with typical frequency of up to 2.5 MHz for
            MII MDC. The input clock, typically provided by HAL, is further
            divided by ENET according to setting of ENET MSCR register in order to
            provide frequency within 2.5 MHz range."
     }

    cdl_option CYGHWR_HAL_FREESCALE_ENET_E0_1588_PORT {
        display "IEEE 1588 Port"
        active_if CYGSEM_DEVS_ETH_FREESCALE_ENET_1588
        parent CYGSEM_DEVS_ETH_FREESCALE_ENET_1588
        flavor data
        default_value { "B" }
        legal_values { "B" "C" "User" }
        description "
            Digital I/O provided by HAL for ENET IEEE 1588 timers."
    }

    cdl_component CYGHWR_DEVS_DISK_FREESCALE_USDHC {
        display "SDHC Disk"
        flavor none

        active_if CYGPKG_DEVS_DISK_FREESCALE_USDHC

    }

    cdl_component CYGHWR_HAL_DEVS_IRQ_PRIO_SCHEME {
        display "Interrupt priority scheme"
        flavor none
        description "Consolidated interrupt priority scheme setting."
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
            Global build options including control over
            compiler flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . CYGBLD_ARCH_CFLAGS .
                            "-Wno-comment -mcpu=cortex-a9 -mfpu=neon -g -O0 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -ffreestanding" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { CYGBLD_ARCH_LDFLAGS . "-mcpu=cortex-a9 -mfpu=neon -static -n -g -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" } 
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image."
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }
}
