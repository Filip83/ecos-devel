# ====================================================================
#
#      uart_ehci_serial.cdl
#
#      eCos serial ehci Freescale Kinetis configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Contributors:   
# Date:           2017-03-28
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_DEVS_EHCI_SERIAL_FREESCALE {
    display       "Freescale uart ehci serial device drivers"

    implements    CYGINT_DEVS_EHCI_KINETIS
    implements    CYGINT_HAL_DMA
    parent		  CYGPKG_IO_EHCI

    requires      CYGPKG_IO_SERIAL_FREESCALE_UART_HDR
    requires      CYGPKG_ERROR
    requires      CYGPKG_HAL_FREESCALE_EDMA
    include_dir   cyg/io
    description   "
           This option enables the ehci serial device drivers for the
           Freescale kinetis uart."
    

    compile       -library=libextras.a   uart_ehci_serial.c

    #define_proc {
    #    puts $::cdl_system_header "/***** serial driver proc output start *****/"
    #     puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_ehci_serial_avr32_uc3c.h>"
    #    puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    #}

    cdl_option CYGDAT_DEVS_EHCI_SERIAL_FREESCALE_NAME {
        display       "Device name for ehci serial driver."
        flavor        data
        default_value {"\"/dev/ehci\""}
        description   "
            This option specifies the name of the ehci serial device."
    }

    cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_BAUD {
        display       "Baud rate for the ehci serial driver."
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 115200
        description   "
            This option specifies the default baud rate (speed) for the 
            ehci driver."
    }

    cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_ISR_PRI {
        display "Interrupt priority"
        flavor        data
        default_value 0x90
        legal_values  { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80 
            0x90  0xA0 0xB0 0xC0 0xD0 0xE0 }
    }

    cdl_component CYGHWR_DEVS_EHCI_SERIAL_FREESCALE_TX_DMA_CHAN {
        display "TX DMA channel"
        flavor data
        default_value 8
        legal_values { 0 to (CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM-1) }
        description "DMA channel assigned to the trasmitter of ehci"

        cdl_component CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_TX_DMA_PRI {
            display "Transmit DMA channel priority"
            flavor data
            legal_values  { 0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 255 }
            default_value 255
            description "
            DMA can work in either round robin or preeptve arbitration
            mode. In preemptive mode, DMA each channel has unique priority,
            lower number meaning lower priority.
            255 is a phony meaning \"default channel priority\"."
        }

        cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_TX_DMA_ECP {
            display "Enable channel preemption"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }

        cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_TX_DMA_DPA {
            display "Disable preempt ability"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }

        cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_TX_DMA_ISR_PRI {
                display "TX DMA channel interrupt priority"
                flavor        data
                default_value 0x90
                legal_values  { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80 
                    0x90  0xA0 0xB0 0xC0 0xD0 0xE0 }
        }
    }

    cdl_component CYGHWR_DEVS_EHCI_SERIAL_FREESCALE_RX_DMA_CHAN {
        display "RX DMA channel"
        flavor data
        default_value 9
        legal_values { 0 to (CYGNUM_HAL_FREESCALE_EDMA_CHAN_NUM-1) }
        description "DMA channel assigned to the receiver of ehci"

        cdl_component CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_RX_DMA_PRI {
            display "Receive DMA channel priority"
            flavor data
            legal_values { 0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 255 }
            default_value 255
            description "
            DMA can work in either round robin or preeptve arbitration
            mode. In preemptive mode, DMA each channel has unique priority,
            lower number meaning lower priority.
            255 is a phony meaning \"default channel priority\"."
        }

        cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_RX_DMA_ECP {
            display "Enable channel preemption"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }

        cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_RX_DMA_DPA {
            display "Disable preempt ability"
            flavor data
            legal_values { 0 1 }
            default_value 0
        }

        cdl_option CYGNUM_DEVS_EHCI_SERIAL_FREESCALE_RX_DMA_ISR_PRI {
                display "RX DMA channel interrupt priority"
                flavor        data
                default_value 0x90
                legal_values  { 0 0x10 0x20 0x30 0x40 0x50 0x60 0x70 0x80 
                    0x90  0xA0 0xB0 0xC0 0xD0 0xE0 }
            }
    }

    cdl_component CYGPKG_DEVS_EHCI_SERIAL_FREESCALE_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_DEVS_EHCI_SERIAL_FREESCALE_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_EHCI_SERIAL_FREESCALE_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF uart_ehci_serial.cdl
