# ====================================================================
#
#      usart_spi_avr32.cdl
#
#      Atmel AVR32UC3C USART SPI driver configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Date:           2013-05-09
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_USART_SPI_AVR32_UC3C {
    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI
    display       "Atmel AVR32UC3C USART SPI driver"
    requires      CYGPKG_HAL_AVR32
    requires      CYGPKG_ERROR
    hardware
    include_dir   cyg/io
    compile       usart_spi_avr32.c
    compile       -library=libextras.a usart_spi_avr32_init.cxx

    cdl_option CYGHWR_DEVS_USART_SPI_AVR32_UC3C_BUS0 {
        display       "Enable support for USART SPI bus 0"
        flavor        bool
        default_value 0
        description   "Enable this option to add support for the USART0 
                       SPI peripheral." 
    }

    cdl_option CYGHWR_DEVS_USART_SPI_AVR32_UC3C_BUS1  {
        display       "Enable support for USART SPI bus 1"
        flavor        bool
        default_value 0
        description   "Enable this option to add support for the USART1 
                       SPI peripheral." 
    }      

    cdl_option CYGHWR_DEVS_USART_SPI_AVR32_UC3C_BUS2 {
        display       "Enable support for USART SPI bus 2"
        flavor        bool
        default_value 0
        description   "Enable this option to add support for the USART2 
                       SPI peripheral." 
    }

    cdl_option CYGHWR_DEVS_USART_SPI_AVR32_UC3C_BUS3  {
        display       "Enable support for USART SPI bus 3"
        flavor        bool
        default_value 0
        description   "Enable this option to add support for the USART3 
                       SPI peripheral." 
    }

    cdl_option CYGHWR_DEVS_USART_SPI_AVR32_UC3C_BUS4  {
        display       "Enable support for USART SPI bus 4"
        flavor        bool
        default_value 0
        description   "Enable this option to add support for the USART4 
                       SPI peripheral." 
    }

    cdl_component CYGPKG_DEVS_USART_SPI_AVR32_UC3C_OPTIONS {
        display "Atmel AVR32 USART SPI driver build options"
        flavor  none
        description   "
	        Package specific build options including control over
	        compiler flags used only in building this package,
	        and details of which tests are built."

        cdl_option CYGPKG_DEVS_USART2_SPI_AVR32_UC3C_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the SPI device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_USART2_SPI_AVR32_UC3C_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the SPI device. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF usart_spi_avr32.cdl
