# ====================================================================
#
#      telnetd.cdl
#
#      TELNETD configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2002 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Mike Jones <mike@proclivis.com>
# Original data:  nickg
# Contributors:   
# Date:           2014-01-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_TELNETD {
    display       "TELNET Daemon"
    parent        CYGPKG_NET
    doc           ref/net-telnetd.html
    include_dir   cyg/telnetd
    requires      CYGPKG_IO
    requires      { 0 != CYGINT_ISO_STDLIB_STRCONV }
    requires      { 0 != CYGINT_ISO_STDIO_FORMATTED_IO }
    requires      { 0 != CYGINT_ISO_STRING_STRFUNCS }
    requires      { 0 != CYGINT_ISO_ERRNO }
    requires      { 0 != CYGINT_ISO_ERRNO_CODES }
    requires      CYGPKG_NET
    description   "
        TELNET Daemon. This is an embedded TELNET server for use with
        applications in eCos. This server is specifically aimed at
        the remote control and monitoring requirements of embedded
        applications. It is NOT intended to be a general purpose server for
        operating a standard shell."

    compile telnetd.cxx
    compile -library=libextras.a init.cxx

    cdl_option CYGNUM_TELNETD_SERVER_PORT {
        display "TELNET port"
        flavor   data
        default_value 23
        description "TELNET port to which browsers will connect.
                     This defaults to the standard port 23, but may
                     be changed to any other port number if required."
    }
    
    cdl_option CYGNUM_TELNETD_THREAD_COUNT {
        display "TELNETD thread count"
        flavor data
        default_value 1
        description "The TELNET server can be configured to use more than
                     one thread to service requests. This is useful if you
                     expect have several simultaneous users. For most purposes, 
                     just one thread is perfectly adequate."
    }

    cdl_option CYGNUM_TELNETD_THREAD_PRIORITY {
        display "THREAD thread priority"
        flavor data
        default_value { CYGNUM_KERNEL_SCHED_PRIORITIES/2 }
        legal_values 0 to CYGNUM_KERNEL_SCHED_PRIORITIES
        description "The THREAD server threads can be run at any priority.
                     The exact priority depends on the importance of the
                     server relative to the rest of the system. The default
                     is to put it in the middle of the priority range to provide
                     reasonable response without impacting genuine high
                     priority threads."
    }

    cdl_option CYGNUM_TELNETD_THREAD_STACK_SIZE {
        display "TELNETD thread stack size"
        flavor data
        default_value 2048
        description "This is the amount of stack to be allocated for each
                     of the TELNETD threads. This quantity is in addition to the values
                     of CYGNUM_HAL_STACK_SIZE_MINIMUM and
                     CYGNUM_TELNETD_SERVER_BUFFER_SIZE."
    }

    cdl_option CYGNUM_TELNETD_SERVER_BUFFER_SIZE {
        display "TELNETD server buffer size"
        flavor data
        default_value 256
        description "This defines the size of the buffer used to receive the first
                     line of each TELNET request. If you expect to use particularly
                     long commands, this should be increased."
    }

    cdl_option CYGNUM_TELNETD_SERVER_AUTO_START {
       display  "Autostart TELNETD"
       default_value 1
       description  "This option causes the TELNET Daemon to be started
                     automatically during system initialization. If this option
                     is not set then the application must start the daemon
                     explicitly by calling cyg_telnetd_startup()."
    }

    cdl_option CYGNUM_TELNETD_SERVER_DELAY {
        display "TELNETD server startup delay"
        flavor data
        default_value 0
        description "This defines the number of system clock ticks that the TELNET
                     server will wait before initializing itself and spawning any
                     extra server threads. This is to give the application a chance
                     to initialize properly without any interference from the TELNETD."
    }
    
    cdl_component CYGPKG_TELNETD_TESTS {
        display "TELNETD tests"
        flavor  data
        no_define
        calculated { 
	    "tests/telnetd1"
        }
        description   "
                This option causes the building of a simple test server."
    }

    cdl_component CYGPKG_TELNETD_COMMANDS {
        display "TELNET server command options"
        flavor  none
	    no_define

        cdl_component CYGPKG_TELNETD_COMMAND_ECHO {
            display "Support the echo command"
            flavor bool
            default_value 1
            description   "
                This option adds an echo command to telnet."
        }

        cdl_component CYGPKG_TELNETD_COMMAND_LUA {
            display "Support Sh Lua"
            flavor bool
            active_if CYGPKG_SH_COMMAND_LUA
            default_value { 0 }
            description   "
                This option adds lua support."                
        }

        cdl_component CYGPKG_TELNETD_COMMAND_DLMALLOC {
            display "Doug Lea Malloc"
            requires (CYGIMP_MEMALLOC_MALLOC_DLMALLOC && \
                CYGIMP_MEMALLOC_ALLOCATOR_DLMALLOC_SAFE_MULTIPLE)
            flavor bool
            default_value { 0 }
            description "
            This option replaces the standard alloc with an instance of 
            dlmalloc that uses its own memory assignment. A dlmalloc
            pool is passed to a shell command and recycled after the command
            completes."
            
             cdl_option CYGPKG_TELNETD_COMMAND_DLMALLOC_SIZE {
                 display "Size of dlmalloc heap"
                 active_if CYGPKG_TELNETD_COMMAND_DLMALLOC
                 flavor data
                 default_value { 10000 }
                 description "
                     Size of memory reserved for a command. Will
                     reserve this size memory for each telnetd
                     thread."
             }
        }

        cdl_component CYGPKG_TELNETD_COMMAND_SH {
            display "Support Sh"
        flavor bool
        active_if CYGPKG_SH
        default_value 0
            description   "
                This option adds sh support."
        }
    }
    
    cdl_component CYGPKG_TELNETD_OPTIONS {
        display "TELNET server build options"
        flavor  none
	no_define

        cdl_option CYGPKG_TELNETD_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the TELNET server package.
	        These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_TELNETD_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the TELNET server package. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF telnetd.cdl
