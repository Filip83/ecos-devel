#==========================================================================
#
#       beep_avr32.cdl
#
#       eCos configuration data for the Atmel AVR32 beeper driver
#
#==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
#==========================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    Filip
# Contributors:
# Date:         2017-04-05
# Purpose:
# Description:  Beeper driver for Frescale Kinetis
#
#####DESCRIPTIONEND####
#
#==========================================================================

cdl_package CYGPKG_DEVS_BEEP_KINETIS {
    display     "Beeper driver."
    requires    CYGPKG_IO
    
    include_dir   cyg/io

    compile       -library=libextras.a beep_kinetis.c

    description "Beeper driver for piezo-electric beeper. This dreiver
                 use Kinetis timer to generate beeper frequncy in wave generation
                 mode. The timer is as well used to generate beeper beep interval"

    cdl_component CYGPKG_DEVS_BEEP_OPTIONS {
        display "options"
        flavor  none
        no_define

        cdl_option CYGPKG_DEVS_BEEP_CFLAGS {
            display       "Additional compiler flags"
            flavor        data
            no_define
            default_value { "" }
            description "
               This option modifies the set of compiler flags for
               building the keypad driver package. These flags
               are used in addition to the set of global flags."
        }
    }

    cdl_option CYGDAT_DEVS_BEEP_NAME {
        display "Device name for the beeper driver"
        flavor data
        default_value {"\"/dev/beep\""}
        description " This option specifies the name of the beeper device"
    }

    cdl_option CYGDAT_DEVS_BEEP_DEFAULT_TIME {
        display "Default beeping timer in ms"
        flavor data
        legal_values     100 to 3000
        default_value { 500 }
    }

    cdl_option CYGDAT_DEVS_BEEP_DEFAULT_FREQUENCY {
        display "Beeper frequncy in Hz"
        flavor data
        legal_values     500 to 10000
        default_value { 4000 }
    }

    cdl_option CYGNUM_DEVS_BEEP_TIMER {
        display "Beeper timer to use FTM0 to FTM2"
        flavor data
        legal_values     0 to 2
        default_value { 0 }
    }

    cdl_option CYGNUM_DEVS_BEEP_CHANNEL {
        display "Timer channel to use"
        flavor data
        legal_values     0 to 7
        default_value { 0 }
    }

    cdl_option CYGNUM_DEVS_BEEP_KINETIS_ISR_PRI {
        display "Interrupt priority"
        flavor data
        calculated 0x90
        description "Interrupt priority is set to defalut value"
    }

    cdl_option CYGDAT_DEVS_BEEP_OUTPUT {
        display "Enable beper driver debug utput"
        flavor data
        legal_values  0 to 3
        default_value { 0 }
    }
}
