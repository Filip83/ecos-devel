# ====================================================================
#
#      nmea_lib.cdl
#
#      NMEA lib configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Contributors:
# Date:           2016-05-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_NMEA_LIB {
    display       "NMEA parser package"
    description   "
                  This package provides support for NMEA
                  messages processing."
    #include_dir   cyg/compress

    requires      CYGPKG_ISOINFRA

    compile       context.c  generate.c  generator.c  gmath.c  info.c  
    compile       parse.c  parser.c  sentence.c  time.c  tok.c

# ====================================================================

  cdl_component CYGPKG_NMEA_LIB_BUFFER_OPTIONS {
      display "NMEA lib package buffers options"
	    flavor  none
	    no_define
	    description   "
		Package parse and time parse buffer size option."
	    
	    
	cdl_option CYGNUM_NMEA_LIB_CONVSTR_BUF_SIZE {
		display       "Sizeof to int converstion buffer in bytes"
		flavor        data
		legal_values  16 to 1024
		default_value 64
		description   "This buffer is allocen on heap
		             and is used in nmea_atoi function."
	    }
	    
	cdl_option CYGNUM_NMEA_LIB_TIMEPARSE_BUF_SIZE {
		display       "Sizeof buffer, in bytes, for time in text form"
		flavor        data
		legal_values  16 to 1024
		default_value 64
		description   "This buffer is allocen on heap
		             and is used to contain time date from NMEA message as text."
	    }
	    
	cdl_option CYGNUM_NMEA_LIB_DEF_PARSEBUFF_SIZE {
	    display       "Sizeof parser buffer"
	    flavor        data
	    legal_values  256 to 10240
	    default_value 1024
	    description   "This buffer is used to fill data in before parsing.
			    This macro is as well used to construct buffers on
			    heap in trace and error messages."
	}
	}

    cdl_component CYGPKG_NMEA_LIB_OPTIONS {
        display "NMEA lib package build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."

        cdl_option CYGPKG_NMEA_LIB_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_NMEA_LIB_LDFLAGS_ADD {
            display "Additional linker flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of linker flags for
                building this package. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_NMEA_LIB_LDFLAGS_REMOVE {
            display "Suppressed linker flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of linker flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }
	
    }

}

# ====================================================================
# EOF nmea_lib.cdl
