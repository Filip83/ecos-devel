# ====================================================================
#
#      ser_freescale_uart.cdl
#
#      eCos serial Freescale UART configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Mike Jones <mike@proclivis.com>
# Contributors:   Ilija Kocho <ilijak@siva.com.mk>
# Original data:
# Contributors:
# Date:           203-08-08
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_FREESCALE_UARTA {
    display       "Freescale UARTA device driver"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    requires      CYGPKG_IO_SERIAL_FREESCALE_UARTA_HDR
    requires      CYGPKG_ERROR

    include_dir   cyg/io

    description   "
        This option enables the serial device drivers for the
        Freescale UART, an on-chip serial controller found on 
        iMX6, etc."

    compile       -library=libextras.a   ser_freescale_uart.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_freescale_uarta.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    # Support up to 5 on-chip UART modules.
    for { set ::channel 0 } { $::channel < 4 } { incr ::channel } {

        cdl_interface CYGINT_IO_SERIAL_FREESCALE_UART[set ::channel] {
            display     "Platform provides UART [set ::channel]"
            flavor      bool
            description "
                This interface will be implemented if the specific
                controller being used has on-chip UART [set ::channel], and if
                that UART is accessible on the target hardware."
        }

        cdl_component CYGPKG_IO_SERIAL_FREESCALE_UART[set ::channel] {
            display       "Freescale UART port [set ::channel] driver"
            flavor        bool
            active_if     CYGINT_IO_SERIAL_FREESCALE_UART[set ::channel]
            default_value CYGINT_IO_SERIAL_FREESCALE_UART[set ::channel]
            implements    CYGINT_IO_SERIAL_TTY_TTY[set ::channel]
            description   "
                This option includes the serial device driver for Freescale
                UART port [set ::channel]."

            cdl_option CYGDAT_IO_SERIAL_FREESCALE_UART[set ::channel]_NAME {
                display       "Device name for Freescale UART port [set ::channel]"
                flavor        data
                default_value [ format {"\"/dev/ser%d\""} $::channel ]
                description   "
                    This option specifies the device name for
                    Freescale UART port [set ::channel]."
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART[set ::channel]_BAUD {
                display       "Baud rate for the Freescale UART port [set ::channel] driver"
                flavor        data
                legal_values  { 300 600 1200 2400 4800 9600 14400 19200 38400
                    57600 115200 230400 }
                default_value 38400
                description "
                    This option specifies the default baud rate for the
                    Freescale UART port [set ::channel]."
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART[set ::channel]_BUFSIZE {
                display       "Buffer size for the Freescale UART port [set ::channel] driver"
                flavor        data
                legal_values  0 to 8192
                default_value 128
                description   "
                    This option specifies the size of the internal buffers used
                    for Freescale UART port [set ::channel]."
            }

            cdl_option CYGNUM_IO_SERIAL_FREESCALE_UART[set ::channel]_INT_PRIORITY {
                display      "Freescale UART port [set ::channel] interrupt priority"
                flavor       data
                default_value CYGNUM_IO_SERIAL_FREESCALE_UART[set ::channel]_INT_PRIORITY_SP
                description   "
                    This option selects the interupt priority for the
                    Freescale UART [set ::channel] interrupts."
            }
        }
    }

    cdl_component CYGDAT_IO_SERIAL_TTY_ADD_INL {
        display "Freescale TTY devices beyond #3"
        parent CYGPKG_IO_SERIAL
        active_if CYGPKG_IO_SERIAL_TTY
        flavor data
        calculated { "<cyg/io/ser_freescale_uart_tty_add.inl>" }


        cdl_component CYGPKG_IO_SERIAL_TTY_TTY4 {
            display       "TTY mode channel #4"
            flavor        bool
            parent        CYGPKG_IO_SERIAL_TTY
            active_if     CYGPKG_IO_SERIAL_TTY
            default_value 0
            description   "
                This option causes '/dev/tty4', which is provided by Freescale
                UART, to be included in the standard drivers."

            cdl_option CYGDAT_IO_SERIAL_TTY_TTY4_DEV {
                display       "TTY mode channel #4 device"
                flavor        data
                default_value { "\"/dev/ser4\"" }
                description   "
                    This option selects the physical device to use for
                    '/dev/tty4'."
            }
        }
    }

    cdl_component CYGDAT_IO_SERIAL_TERMIOS_ADD_INL {
        display "Freescale TERMIOS devices beyond #3"
        parent CYGPKG_IO_SERIAL
        active_if CYGPKG_IO_SERIAL_TERMIOS
        flavor data
        calculated { "<cyg/io/ser_freescale_uart_termiostty_add.inl>" }

        cdl_component CYGPKG_IO_SERIAL_TERMIOS_TERMIOS4 {
            display       "Termios TTY channel #4"
            flavor        bool
            default_value 0
            implements    CYGINT_IO_SERIAL_TERMIOS_TERMIOS_TTY
            parent        CYGPKG_IO_SERIAL_TERMIOS
            active_if     CYGPKG_IO_SERIAL_TERMIOS
            description   "
                This option causes '/dev/termios4' to be included in the
                standard drivers."

            cdl_option CYGDAT_IO_SERIAL_TERMIOS_TERMIOS4_DEV {
                display       "Termios TTY channel #4 device"
                flavor        data
                default_value {"\"/dev/ser4\""}
                description   "
                    This option selects the physical device to use for
                    '/dev/termios4'."
            }
        }

    }

    cdl_component CYGPKG_IO_SERIAL_FREESCALE_UART_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
            Package specific build options including control over
            compiler flags used only in building this package,
            and details of which tests are built."

        cdl_option CYGPKG_IO_SERIAL_FREESCALE_UART_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are
                used in addition to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_FREESCALE_UART_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are
                removed from the set of global flags if present."
        }
    }
}

# EOF ser_freescale_uart.cdl
