# ====================================================================
#
#      adc_avr32.cdl
#
#      eCos AVR32UC3C ADC configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2008 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Contributors:
# Date:           2012-11-15
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_DEVS_ADC_AVR32_UC3C {
    display     "ADC hardware device driver for AVR32 family of controllers"

    parent      CYGPKG_IO_ADC
    active_if   CYGPKG_HAL_AVR32
    description "
           This package provides a generic ADC device driver for the on-chip
           ADC peripherals in AVR32UC3C processors."

    include_dir cyg/io
    compile     -library=libextras.a adc_uc3c.c

    define_proc {
      puts $::cdl_system_header "#define CYGDAT_DEVS_ADC_AVR32_UC3C_INL <cyg/io/adc_uc3c.inl>"
    }

    #
    # Primary ADC ( ADC0 )
    #
    cdl_component CYGPKG_DEVS_ADC_AVR32_UC3C_ADC0 {
        display       "Atmel AVR32 ADC port 0 driver"
        flavor        bool
        default_value 1
        description "
           This option includes the device driver for the on-chip ADC 0 of the
           AVR32UC3C processors. For now only one sequncer is implemented e.g.
           only ADCIN0 to ADCIN7 can be used and non diferencial inputs."


        cdl_interface CYGINT_DEVS_ADC_AVR32_UC3C_ADC0_CHANNELS {
          display "Number of ADC0 channels"
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_PRESCAL {
            display       "ADC clock prescaller setting"
            flavor        data
            legal_values  0 to 512
            default_value 128
            description   "
               This option sets the AVR32UC3C ADC PRESCAL value.
               ADCClock = MCK / ((PRESCAL + 1) * 2)"
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_STARTUP_TIME {
            display       "ADC start-up time"
            flavor        data
            legal_values  0 to 64
            default_value 0
            description   "
               This option sets the AVR32UC3C ADC start-up time value.
               ADC start-up time = (STARTUP+1) * 32 / ADCClock"
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_MUX_SETTLE_TIME {
            display       "ADC mux settle time 1.5"
            flavor        bool
            default_value 0
            description   "
               This option sets the AVR32UC3C ADC muxes settle time."
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_EXTERNAL_REFERENCE {
            display       "Forece use external refernce ADCRERFN/P"
            flavor        bool
            default_value 0
            description   "
               This option foce the AVR32UC3C ADC to use external
               reference on ADCREFN and ADCREFP pads."
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_REFERENCE {
            display       "ADC reference select"
            active_if     !CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_EXTERNAL_REFERENCE
            flavor        data
            legal_values  {"INT1V" "INT0_6VDDANA" "EXTADCERF0" "EXTADCREF1"}
            default_value { "INT0_6VDDANA"}
            description   "
               This options select the ADC reference."
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_SAH_DISABLE {
            display       "Disable sample and hold"
            flavor        bool
            default_value 0
            description   "
               When this option is enabled the internal smple and
               hold circuit is disabled as well as sequencer 1.
               The adc latency is decreased by one ADC clock."
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_SIGNLE_SEQUENCER_ENABLE {
            display       "Enable single sequncer mode"
            flavor        bool
            default_value 0
            description   "
               When this option enable single sequencer mode to increase
               the number of conversion per sequence."
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_SLEEP_DISABLE {
            display       "Disable sleep mode"
            flavor        bool
            default_value 0
            description   "
               This option disable sllep mode betwen conversions."
        }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_INTPRIO {
            display       "Interrupt priority"
            flavor        data
            legal_values  0 to 3
            default_value 0
       }

        cdl_option CYGNUM_DEVS_ADC_AVR32_UC3C_ADC0_DEFAULT_RATE {
            display "Default sample rate"
            flavor   data
            legal_values 0 to 131072
            default_value 100
            description "
               The driver will be initialized with the default sample rate.
               If you raise the default sample rate you might need to increase
               the buffer size for each channel. If sample rate is zero the sample
               is taken only after new setting of sampling rate to zero or
               by setiing any higher number the sample gnerator is neabled."
        }

        # Support up to 8 ADC channels
        for { set ::channel 0 } { $::channel < 8 } { incr ::channel } {

            cdl_component CYGPKG_DEVS_ADC_AVR32_UC3C_ADC0_CHANNEL[set ::channel] {
                display        "Access ADC channel [set ::channel]"
                flavor          bool
                default_value   [set ::channel] == 0
                implements      CYGINT_DEVS_ADC_AVR32_UC3C_ADC0_CHANNELS
                description "
                   If the application needs to access the on-chip ADC
                   channel [set ::channel] via an eCos ADC driver then
                   this option should be enabled."

                cdl_option CYGDAT_DEVS_ADC_AVR32_UC3C_ADC0_CHANNEL[set ::channel]_NAME {
                    display "Device name"
                    flavor      data
                    default_value   [format {"\"/dev/adc0%d\""} $::channel]
                    description "
                       This option controls the name that an eCos application
                       should use to access this device via cyg_io_lookup(),
                       open(), or similar calls."
                }

                cdl_option CYGDAT_DEVS_ADC_AVR32_UC3C_ADC0_CHANNEL[set ::channel]_BUFSIZE {
                    display "Size of data buffer"
                    flavor  data
                    legal_values  0x01 to 0x2000000
                    default_value 16
                    description "
                       This option controls the number of samples the
                       buffer can store. The required RAM depends on the
                       sample size and on the number of samples. If the
                       sample size is <= 8 bit the the required RAM =
                       size of data buffer. If the sample size is 9 or 10
                       bit then required RAM = size of data buffer * 2."
                }
            }
        }
    }

    cdl_option CYGPKG_DEVS_ADC_AVR32_UC3C_DEBUG_LEVEL {
        display "Driver debug output level"
        flavor  data
        legal_values {0 1}
        default_value 0
        description   "
             This option specifies the level of debug data output by
             the AVR32UC3C ADC device driver. A value of 0 signifies
             no debug data output; 1 signifies normal debug data
             output. If an overrun occurred then this can only be
             detected by debug output messages."
    }
}
