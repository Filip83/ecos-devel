# ====================================================================
#
#      kinetis_gpio.cdl
#
#      eCos Frescale Kinetis GPIO configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2008 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Contributors:
# Date:           2019-03-26
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_DEVS_GPIO_KINETIS {
    display     "GPIO hardware device driver for kinetis family of controllers"
    implements  CYGHWR_DEVS_GPIO_KINETIS
    parent      CYGPKG_IO_GPIO
    description "
           This package provides a generic and simple GPIO device driver for the on-chip
           GPIO, PWM, ADC and DAC peripherals in kinetis processors."

    include_dir cyg/io/gpio
    compile     -library=libextras.a   \
	             analogin_api.c		   \
				 analogout_api.c	   \
				 gpio_api.c            \
				 PeripheralPins.c      \
				 port_api.c            \
				 pwmout_api.c

}
