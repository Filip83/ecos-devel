# ====================================================================
#
#      usbs_kinetis.cdl
#
#      USB device driver for the Freescale Kinetis family of processors.
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2006, 2010 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later
## version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License
## along with eCos; if not, write to the Free Software Foundation, Inc.,
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
##
## As a special exception, if other files instantiate templates or use
## macros or inline functions from this file, or you compile this file
## and link it with other works to produce a work based on this file,
## this file does not by itself cause the resulting work to be covered by
## the GNU General Public License. However the source code for this file
## must still be made available in accordance with section (3) of the GNU
## General Public License v2.
##
## This exception does not invalidate any other reasons why a work based
## on this file might be covered by the GNU General Public License.
## -------------------------------------------
## ####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Contributors:
# Date:           2017-04-20
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_DEVS_USB_KINETIS {
    display     "Freescale Kinetis USB Device Driver"
    include_dir "cyg/io/usb"
    parent      CYGPKG_IO_USB
    implements  CYGHWR_IO_USB_SLAVE


    description "
        This package provides a suitable eCos device driver
        for Freescale Kinetis USB.
        The Driver needs 48MHz plus minus 0.25%.
        Buffers are allocated only in the higher level. There
        is no need to configure the endpoints in this CDL, because
        they will be configured dynamical at the set_configuration
        call from the host...
        The endpoints 1..3 can be configured as bulk or interrupt
        IN or OUT endpoint."
        
    cdl_component CYGFUN_DEVS_USB_KINETIS_STLIB_SUPPORT {
        display       "Enable StLib USB messages"
        flavor        bool
        default_value 0

        description   "
            Enable support for StLib to send messages
            about USB state change."
    }
    
    cdl_component CYGFUN_DEVS_USB_KINETIS_EP0 {
        display       "Support the control endpoint 0"
        flavor        bool
        default_value CYGINT_IO_USB_SLAVE_CLIENTS
        requires      CYGPKG_IO_USB CYGPKG_IO_USB_SLAVE

        implements CYGHWR_IO_USB_SLAVE_OUT_ENDPOINTS
        implements CYGHWR_IO_USB_SLAVE_IN_ENDPOINTS

        compile       -library=libextras.a usbc_kinetis.c usbs_kinetis_data.cxx

        description   "
            Enable support for endpoint 0. If this support is disabled
            then the entire USB port is unusable."

    }

    cdl_component CYGPKG_DEVS_USB_KINETIS_DEVTAB_ENTRIES {
        display       "Provide a devtab entry for endpoints"
        active_if     CYGFUN_DEVS_USB_KINETIS_EP0
        default_value 0
        description "
             This component controls if /dev/usb entries will be created."

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP0_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 0"
            flavor        bool
            default_value 0
            requires      CYGPKG_IO
            description "
               If endpoint 0 will only be accessed via the low-level
               USB-specific calls then there is no need for an entry
               in the device table, saving some memory. If the
               application intends to access the endpoint by means
               of open and ioctl calls then a devtab entry is needed."
        }

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP1_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 1"
            flavor        bool
            default_value 1
            requires      CYGPKG_IO
            description "
                If this endpoint will only be accessed via the low-level
                USB-specific calls then there is no need for an entry
                in the device table, saving some memory. If the
                application intends to access the endpoint by means
                of open and read calls then a devtab entry is needed."
        }

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP2_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 2"
            flavor        bool
            default_value 1
            requires      CYGPKG_IO
            description "
                If this endpoint will only be accessed via the low-level
                USB-specific calls then there is no need for an entry
                in the device table, saving some memory. If the
                application intends to access the endpoint by means
                of open and read calls then a devtab entry is needed."


        }

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP3_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 3"
            flavor        bool
            default_value 1
            requires      CYGPKG_IO
            description "
                If this endpoint will only be accessed via the low-level
                USB-specific calls then there is no need for an entry
                in the device table, saving some memory. If the
                application intends to access the endpoint by means
                of open and read calls then a devtab entry is needed."
        }

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP4_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 4"
            flavor        bool
            default_value 0
            requires      CYGPKG_IO
            description "
                If this endpoint will only be accessed via the low-level
                USB-specific calls then there is no need for an entry
                in the device table, saving some memory. If the
                application intends to access the endpoint by means
                of open and read calls then a devtab entry is needed."
        }

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP5_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 5"
            flavor        bool
            default_value 0
            requires      CYGPKG_IO
            description "
                If this endpoint will only be accessed via the low-level
                USB-specific calls then there is no need for an entry
                in the device table, saving some memory. If the
                application intends to access the endpoint by means
                of open and read calls then a devtab entry is needed."
        }

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP6_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 6"
            flavor        bool
            default_value 0
            requires      CYGPKG_IO
            description "
                If this endpoint will only be accessed via the low-level
                USB-specific calls then there is no need for an entry
                in the device table, saving some memory. If the
                application intends to access the endpoint by means
                of open and read calls then a devtab entry is needed."
        }

        cdl_option CYGVAR_DEVS_USB_KINETIS_EP7_DEVTAB_ENTRY {
            display       "Provide a devtab entry for endpoint 7"
            flavor        bool
            default_value 0
            requires      CYGPKG_IO
            description "
                If this endpoint will only be accessed via the low-level
                USB-specific calls then there is no need for an entry
                in the device table, saving some memory. If the
                application intends to access the endpoint by means
                of open and read calls then a devtab entry is needed."
        }


        cdl_option CYGDAT_DEVS_USB_KINETIS_DEVTAB_BASENAME {
            display       "Base name for devtab entries"
            flavor        data
            default_value { "\"/dev/usbs\"" }
            description "
                If the Kinetis USB device driver package provides devtab
                entries for any of the endpoints then this option gives
                control over the names of these entries. By default the
                endpoints will be called \"/dev/usbs0c\", \"/dev/usbs3w\"
                and \"/dev/usbs4r\" (assuming all three endpoints are
                enabled. The common part \"/dev/usbs\" is determined
                by this configuration option. It may be necessary to
                change this if there are multiple USB slave-side
                devices on the target hardware to prevent a name clash."
        }
    }
}
