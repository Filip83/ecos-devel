# ====================================================================
#
#      fb_st7565.cdl
#
#      Framebuffer device driver for the ST7565 target.
#
# ====================================================================
# ####ECOSGPLCOPYRIGHTBEGIN####                                             
# -------------------------------------------                               
# This file is part of eCos, the Embedded Configurable Operating System.    
# Copyright (C) 2008, 2009 Free Software Foundation, Inc.                         
#
# eCos is free software; you can redistribute it and/or modify it under     
# the terms of the GNU General Public License as published by the Free      
# Software Foundation; either version 2 or (at your option) any later       
# version.                                                                  
#
# eCos is distributed in the hope that it will be useful, but WITHOUT       
# ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or     
# FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License     
# for more details.                                                         
#
# You should have received a copy of the GNU General Public License         
# along with eCos; if not, write to the Free Software Foundation, Inc.,     
# 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.             
#
# As a special exception, if other files instantiate templates or use       
# macros or inline functions from this file, or you compile this file       
# and link it with other works to produce a work based on this file,        
# this file does not by itself cause the resulting work to be covered by    
# the GNU General Public License. However the source code for this file     
# must still be made available in accordance with section (3) of the GNU    
# General Public License v2.                                                
#
# This exception does not invalidate any other reasons why a work based     
# on this file might be covered by the GNU General Public License.          
# -------------------------------------------                               
# ####ECOSGPLCOPYRIGHTEND####                                               
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):     Filip  <filip.gnu@gmail.com>
# Date:          2016-11-24
#
#####DESCRIPTIONEND####
#========================================================================

cdl_package CYGPKG_DEVS_FRAMEBUF_ST7565 {
    display		"ST7565 Target Framebuffer device driver"
    parent		CYGPKG_IO_FRAMEBUF
    active_if		CYGPKG_IO_FRAMEBUF
    implements		CYGINT_IO_FRAMEBUF_DEVICES
    implements		CYGHWR_IO_FRAMEBUF_FUNCTIONALITY_DOUBLE_BUFFER
    hardware
    include_dir         cyg/io
    
    compile       -library=libextras.a fb_st7565.c
    description "
        This package provides a framebuffer device driver for the
        ST7565 target."

    cdl_option CYGNUM_DEVS_FRAMEBUF_ST7565_FB_WIDTH {
        display		"Display width"
        flavor 		data
        default_value	132
        legal_values	16 to 132
    }

    cdl_option CYGNUM_DEVS_FRAMEBUF_ST7565_FB_HEIGHT {
        display		"Display height"
        flavor 		data
        default_value	32
        legal_values	8 to 64
    }

    cdl_option CYGNUM_DEVS_FRAMEBUF_ST7565_FB_STRIDE {
        display		"Display stride"
        flavor 		data
        default_value	4
        legal_values	1 to 4
        description "This value respond to nuber of visible display pages."
    }
    
    cdl_option CYGNUM_DEVS_FRAMEBUF_ST7565_FB_ENDIAN {
        display		"Display endian"
        flavor 		data
        default_value	"CYG_FB_FLAGS0_LE"
        legal_values	"CYG_FB_FLAGS0_LE"
        description "This option cannot be modified by user."
    }

    cdl_option CYGNUM_DEVS_FRAMEBUF_ST7565_ENABLE_BACKLIGHT_CONTROL {
        display		"Enable driver to control back light"
        flavor 		bool
        default_value	1
    }

    cdl_option CYGNUM_DEVS_FRAMEBUF_ST7565_BACKLIGHT_PIN {
        display		"Pin name used to control backlight"
        flavor 		data
        default_value	"AVR32_PIN_PC15"
        active_if       CYGNUM_DEVS_FRAMEBUF_ST7565_ENABLE_BACKLIGHT_CONTROL
    }

    cdl_option CYGNUM_DEVS_FRAMEBUF_ST7565_A0_PIN {
        display		"Display pin to control command/data"
        flavor 		data
        default_value	"AVR32_PIN_PC15"
    }

    cdl_component CYGPKG_DEVS_FRAMEBUF_ST7565_OPTIONS {
        display "Framebuffer build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building the synthetic
            target framebuffer device driver."

        cdl_option CYGPKG_DEVS_FRAMEBUF_ST7565_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for building
                the synthetic target framebuffer device driver. These flags
                are used in addition to the set of global flags."
        }

        cdl_option CYGPKG_DEVS_FRAMEBUF_ST7565_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for building
                the synthetic target framebuffer device driver. These flags
                are removed from the set of global flags if present."
        }
    }
}