# ====================================================================
#
#      ser_ar32.cdl
#
#      eCos serial Atmel AVR32UC3C configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Filip
# Contributors:   
# Date:           2016-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_EHCI_SERIAL_AVR32_UC3C {
    display       "Atmel AVR32UC3C ehci serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_AVR32

    requires      CYGPKG_ERROR
    include_dir   cyg/io
    description   "
           This option enables the ehci serial device drivers for the
           Atmel AVR32."
    

    compile       -library=libextras.a   avr32_ehci_serial.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_ehci_serial_avr32_uc3c.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_EHCI_SERIAL_AVR32_SERIAL0 {
    display       "Atmel AVR32UC3C0512 serial port 0 driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for the Atmel AVR32 
        port 0."


    cdl_option CYGDAT_IO_EHCI_SERIAL_AVR32_SERIAL0_NAME {
        display       "Device name for Atmel AVR32UC3C serial port 0 driver"
        flavor        data
        default_value {"\"/dev/ehci0\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AVR32UC3C port 0."
    }

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL0_BAUD {
        display       "Baud rate for the Atmel AVR32UC3C serial port 0 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the 
            Atmel AVR32UC3C port 0."
    }

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL0_FLOW_CONTROL {
        display       "Enable serial flow contrl RTS CTS on serial port 0"
        flavor        bool
        default_value 0
        description   "
            Enable hardware flow control for serial port."

       implements    CYGINT_IO_EHCI_SERIAL_FLOW_CONTROL_HW
       
    }
}

cdl_component CYGPKG_IO_EHCI_SERIAL_AVR32_SERIAL1 {
    display       "Atmel AVR32UC3C serial port 1 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the Atmel AVR32UC3C 
        port 1 (serial B)."


    cdl_option CYGDAT_IO_EHCI_SERIAL_AVR32_SERIAL1_NAME {
        display       "Device name for Atmel AVR32UC3C serial port 1 driver"
        flavor        data
        default_value {"\"/dev/ehci1\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AVR32UC3C port 1."
    }

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL1_BAUD {
        display       "Baud rate for the Atmel AVR32UC3C serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            Atmel AVR32UC3C port 1."
    }


    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL1_FLOW_CONTROL {
        display       "Enable serial flow contrl RTS CTS on serial port 1"
        flavor        bool
        default_value 0
        description   "
            Enable hardware flow control for serial port."

       implements    CYGINT_IO_EHCI_SERIAL_FLOW_CONTROL_HW
       
    }
}

cdl_component CYGPKG_IO_EHCI_SERIAL_AVR32_SERIAL2 {
    display       "Atmel AVR32UC3C serial port 2 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the Atmel AVR32UC3C 
        port 2 (serial C)."

    cdl_option CYGDAT_IO_EHCI_SERIAL_AVR32_SERIAL2_NAME {
        display       "Device name for Atmel AVR32UC3C serial port 1 driver"
        flavor        data
        default_value {"\"/dev/ehci2\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AVR32UC3C port 2."
    }

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL2_BAUD {
        display       "Baud rate for the Atmel AVR32UC3C serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            Atmel AVR32UC3C port 2."
    }
    

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL2_FLOW_CONTROL {
        display       "Enable serial flow contrl RTS CTS on serial port 2"
        flavor        bool
        default_value 0
        description   "
            Enable hardware flow control for serial port."

       implements    CYGINT_IO_EHCI_SERIAL_FLOW_CONTROL_HW
       
    }
}

cdl_component CYGPKG_IO_EHCI_SERIAL_AVR32_SERIAL3 {
    display       "Atmel AVR32UC3C serial port 3 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the Atmel AVR32UC3C 
        port 2 (serial C)."

    cdl_option CYGDAT_IO_EHCI_SERIAL_AVR32_SERIAL3_NAME {
        display       "Device name for Atmel AVR32UC3C serial port 1 driver"
        flavor        data
        default_value {"\"/dev/ehci3\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AVR32UC3C port 2."
    }

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL3_BAUD {
        display       "Baud rate for the Atmel AVR32UC3C serial port 1 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            Atmel AVR32UC3C port 2."
    }

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL3_FLOW_CONTROL {
        display       "Enable serial flow contrl RTS CTS on serial port 3"
        flavor        bool
        default_value 0
        description   "
            Enable hardware flow control for serial port."

       implements    CYGINT_IO_EHCI_SERIAL_FLOW_CONTROL_HW
       
    }
}

cdl_component CYGPKG_IO_EHCI_SERIAL_AVR32_SERIAL4 {
    display       "Atmel AVR32UC3C serial port 4 driver"
    flavor        bool
    default_value 1
    description   "
        This option includes the serial device driver for the Atmel AVR32UC3C 
        port 2 (serial C)."


    cdl_option CYGDAT_IO_EHCI_SERIAL_AVR32_SERIAL4_NAME {
        display       "Device name for Atmel AVR32UC3C serial port 4 driver"
        flavor        data
        default_value {"\"/dev/ehci\""}
        description   "
            This option specifies the name of the serial device for the 
            Atmel AVR32UC3C port 2."
    }

    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL4_BAUD {
        display       "Baud rate for the Atmel AVR32UC3C serial port 4 driver"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 38400
        description   "
            This option specifies the default baud rate (speed) for the
            Atmel AVR32UC3C port 2."
    }
    
    cdl_option CYGNUM_IO_EHCI_SERIAL_AVR32_SERIAL4_FLOW_CONTROL {
        display       "Enable serial flow contrl RTS CTS on serial port 4"
        flavor        bool
        default_value 0
        description   "
            Enable hardware flow control for serial port."

       implements    CYGINT_IO_EHCI_SERIAL_FLOW_CONTROL_HW
       
    }
    
}

    cdl_component CYGPKG_IO_EHCI_SERIAL_AVR32_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_IO_EHCI_SERIAL_AVR32_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_EHCI_SERIAL_AVR32_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }
}

# EOF avr32_ehci_serial.cdl
