##==========================================================================
##
##      io_gpio.cdl
##
##      Generic GPIO driver layer
##
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
#######DESCRIPTIONBEGIN####
##
## Author(s):    Filp
## Date:         2019-03-26
## Description:  Implements generic layer of GPIO drivers.
##
######DESCRIPTIONEND####
##
##========================================================================*/


cdl_package CYGPKG_IO_GPIO {
    display       "GPIO device drivers"
    parent        CYGPKG_IO
    active_if     CYGPKG_IO
    requires      CYGPKG_ERROR
    include_dir   cyg/io/gpio
    description   "
        This option enables drivers for basic GPIO control. 
		Those drivers are taken from embed OS. This package 
		contains a simple driver for input and output pins,
		ports, PWM and analog in/out. The drivers are 
		implemented as C++ classes. For more details
		see embed OS."

    compile       -library=libextras.a mbed_gpio.c          \
	                                   mbed_pinmap_common.c \
									   BusIn.cpp	        \
									   BusInOut.cpp         \
									   BusOut.cpp
	                       

    cdl_component CYGPKG_IO_GPIO_PORT_DEVICES {
        display       "Enable port device drivers"
        flavor        bool
        default_value 0
        description   "
            This option enables the hardware device drivers
	    for the current platform."

		cdl_component CYGPKG_IO_GPIO_PORT_DEVICES_OUT {
			display       "Enable port out device drivers"
			flavor        bool
			default_value 0
			description   "
				This option enables the hardware device drivers
			for the current platform."
		}

		cdl_component CYGPKG_IO_GPIO_PORT_DEVICES_IN {
			display       "Enable port in device drivers"
			flavor        bool
			default_value 0
			description   "
				This option enables the hardware device drivers
			for the current platform."
		}

		cdl_component CYGPKG_IO_GPIO_PORT_DEVICES_IN_OUT {
			display       "Enable port in/out device drivers"
			flavor        bool
			default_value 0
			description   "
				This option enables the hardware device drivers
			for the current platform."
		}
	}

	cdl_component CYGPKG_IO_GPIO_PWM {
		display       "Enable gpio pwm device drivers"
		flavor        bool
		default_value 0
		description   "
			This option enables the hardware device drivers
		for the current platform."
	}

	cdl_component CYGPKG_IO_GPIO_ANALOG_OUT {
		display       "Enable gpio analog out device drivers"
		flavor        bool
		default_value 0
		description   "
			This option enables the hardware device drivers
		for the current platform."
	}

	cdl_component CYGPKG_IO_GPIO_ANALOG_IN {
		display       "Enable gpio analog in device drivers"
		flavor        bool
		default_value 0
		description   "
			This option enables the hardware device drivers
		for the current platform."
	}
}    
